CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files (x86)\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
20
7 Ground~
168 346 378 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5130 0 0
2
45247.3 0
0
13 Logic Switch~
5 337 232 0 1 11
0 22
0
0 0 21104 0
2 0V
-6 -16 8 -8
2 S1
-26 -7 -12 1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
45247.3 0
0
13 Logic Switch~
5 82 319 0 1 11
0 21
0
0 0 21104 0
2 0V
-6 -16 8 -8
2 B4
-30 -3 -16 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
45247.3 3
0
13 Logic Switch~
5 82 345 0 1 11
0 18
0
0 0 21104 0
2 0V
-6 -16 8 -8
2 B3
-30 -3 -16 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
45247.3 2
0
13 Logic Switch~
5 81 373 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21104 0
2 5V
-6 -16 8 -8
2 B2
-30 -3 -16 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
45247.3 1
0
13 Logic Switch~
5 82 403 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21104 0
2 5V
-6 -16 8 -8
2 B1
-30 -3 -16 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
45247.3 0
0
13 Logic Switch~
5 82 269 0 1 11
0 14
0
0 0 21104 0
2 0V
-6 -16 8 -8
2 A1
-30 -3 -16 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8901 0 0
2
45247.3 0
0
13 Logic Switch~
5 81 239 0 1 11
0 16
0
0 0 21104 0
2 0V
-6 -16 8 -8
2 A2
-30 -3 -16 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7361 0 0
2
45247.3 0
0
13 Logic Switch~
5 82 211 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21104 0
2 5V
-6 -16 8 -8
2 A3
-30 -3 -16 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4747 0 0
2
45247.3 0
0
13 Logic Switch~
5 82 185 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21104 0
2 5V
-6 -16 8 -8
2 A4
-30 -3 -16 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
972 0 0
2
45247.3 0
0
12 Hex Display~
7 532 259 0 16 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3472 0 0
2
45247.3 0
0
5 4071~
219 180 108 0 3 22
0 20 21 9
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
9998 0 0
2
45247.3 0
0
5 4071~
219 181 153 0 3 22
0 19 18 8
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
3536 0 0
2
45247.3 0
0
5 4071~
219 180 199 0 3 22
0 16 17 7
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
4597 0 0
2
45247.3 0
0
5 4071~
219 179 243 0 3 22
0 14 15 6
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
3835 0 0
2
45247.3 0
0
5 4081~
219 183 422 0 3 22
0 14 15 10
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
3670 0 0
2
45247.3 0
0
5 4081~
219 184 382 0 3 22
0 16 17 11
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
5616 0 0
2
45247.3 0
0
5 4081~
219 184 340 0 3 22
0 19 18 12
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
9323 0 0
2
45247.3 0
0
5 4081~
219 185 292 0 3 22
0 20 21 13
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
317 0 0
2
45247.3 0
0
7 74LS157
122 387 323 0 14 29
0 22 13 9 12 8 11 7 10 6
23 5 4 3 2
0
0 0 4848 0
6 74F157
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 0 0 0 0
1 U
3108 0 0
2
45247.3 0
0
31
1 0 0 0 0 0 0 1 0 0 31 3
346 372
349 370
349 368
14 1 2 0 0 4224 0 20 11 0 0 3
419 359
541 359
541 283
13 2 3 0 0 4224 0 20 11 0 0 3
419 341
535 341
535 283
12 3 4 0 0 4224 0 20 11 0 0 3
419 323
529 323
529 283
11 4 5 0 0 4224 0 20 11 0 0 3
419 305
523 305
523 283
3 9 6 0 0 8320 0 15 20 0 0 4
212 243
321 243
321 359
355 359
3 7 7 0 0 4224 0 14 20 0 0 6
213 199
365 199
365 258
326 258
326 341
355 341
3 5 8 0 0 4224 0 13 20 0 0 6
214 153
360 153
360 263
331 263
331 323
355 323
3 3 9 0 0 8320 0 12 20 0 0 6
213 108
355 108
355 268
336 268
336 305
355 305
3 8 10 0 0 4224 0 16 20 0 0 4
204 422
326 422
326 350
355 350
3 6 11 0 0 4224 0 17 20 0 0 4
205 382
332 382
332 332
355 332
3 4 12 0 0 4224 0 18 20 0 0 4
205 340
341 340
341 314
355 314
3 2 13 0 0 4224 0 19 20 0 0 4
206 292
341 292
341 296
355 296
0 1 14 0 0 4096 0 0 15 22 0 3
132 269
132 234
166 234
0 2 15 0 0 4224 0 0 15 23 0 3
117 403
117 252
166 252
0 1 16 0 0 4096 0 0 14 25 0 3
135 239
135 190
167 190
0 2 17 0 0 4224 0 0 14 24 0 3
126 373
126 208
167 208
0 2 18 0 0 4224 0 0 13 26 0 3
121 345
121 162
168 162
0 1 19 0 0 4112 0 0 13 27 0 3
128 211
128 144
168 144
0 1 20 0 0 4096 0 0 12 29 0 3
105 185
105 99
167 99
0 2 21 0 0 4224 0 0 12 28 0 3
113 319
113 117
167 117
1 1 14 0 0 8320 0 7 16 0 0 4
94 269
136 269
136 413
159 413
1 2 15 0 0 0 0 6 16 0 0 4
94 403
126 403
126 431
159 431
1 2 17 0 0 0 0 5 17 0 0 4
93 373
139 373
139 391
160 391
1 1 16 0 0 8320 0 8 17 0 0 4
93 239
142 239
142 373
160 373
1 2 18 0 0 0 0 4 18 0 0 4
94 345
152 345
152 349
160 349
1 1 19 0 0 8320 0 9 18 0 0 4
94 211
147 211
147 331
160 331
1 2 21 0 0 0 0 3 19 0 0 4
94 319
153 319
153 301
161 301
1 1 20 0 0 8320 0 10 19 0 0 4
94 185
153 185
153 283
161 283
1 1 22 0 0 4224 0 2 20 0 0 3
349 232
349 287
355 287
10 0 23 0 0 4224 0 20 0 0 0 2
349 368
345 368
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
