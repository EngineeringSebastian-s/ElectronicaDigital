CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 1
20 Package,Description,
48 C:\Program Files (x86)\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 168 226 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-33 0 -19 8
2 V4
-34 -11 -20 -3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6435 0 0
2
45226.3 1
0
13 Logic Switch~
5 160 365 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-33 0 -19 8
2 V3
-34 -11 -20 -3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5283 0 0
2
45226.3 0
0
13 Logic Switch~
5 167 198 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-33 0 -19 8
2 V2
-34 -11 -20 -3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6874 0 0
2
45226.3 0
0
13 Logic Switch~
5 166 171 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-33 0 -19 8
2 V1
-34 -11 -20 -3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5305 0 0
2
45226.3 0
0
7 Ground~
168 357 296 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
34 0 0
2
45226.3 0
0
5 4049~
219 552 268 0 2 22
0 11 4
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 2 0
1 U
969 0 0
2
45226.3 0
0
5 4049~
219 519 240 0 2 22
0 10 5
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 2 0
1 U
8402 0 0
2
45226.3 0
0
5 4049~
219 466 194 0 2 22
0 9 6
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 2 0
1 U
3751 0 0
2
45226.3 0
0
5 4049~
219 553 169 0 2 22
0 8 7
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 2 0
1 U
4292 0 0
2
45226.3 0
0
8 4-In OR~
219 620 213 0 5 22
0 7 6 5 4 12
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 1 0
1 U
6118 0 0
2
45226.3 0
0
14 Logic Display~
6 701 138 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
34 0 0
2
45226.3 0
0
7 74LS138
19 388 218 0 14 29
0 15 14 13 3 2 2 8 16 17
9 10 18 11 19
0
0 0 5104 0
6 74F138
-21 -61 21 -53
2 U1
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 512 0 0 0 0
1 U
6357 0 0
2
45226.3 0
0
15
6 1 2 0 0 8320 0 12 5 0 0 5
350 254
351 254
351 282
357 282
357 290
5 6 2 0 0 0 0 12 12 0 0 2
350 245
350 254
1 4 3 0 0 4240 0 2 12 0 0 4
172 365
342 365
342 236
356 236
2 4 4 0 0 8320 0 6 10 0 0 4
573 268
595 268
595 227
603 227
2 3 5 0 0 4224 0 7 10 0 0 4
540 240
590 240
590 218
603 218
2 2 6 0 0 4224 0 8 10 0 0 4
487 194
580 194
580 209
603 209
2 1 7 0 0 8320 0 9 10 0 0 4
574 169
595 169
595 200
603 200
7 1 8 0 0 12416 0 12 9 0 0 4
426 191
432 191
432 169
538 169
10 1 9 0 0 4224 0 12 8 0 0 3
426 218
451 218
451 194
11 1 10 0 0 12416 0 12 7 0 0 4
426 227
441 227
441 240
504 240
13 1 11 0 0 12416 0 12 6 0 0 4
426 245
441 245
441 268
537 268
5 1 12 0 0 4224 0 10 11 0 0 3
653 213
653 156
701 156
1 3 13 0 0 4224 0 1 12 0 0 4
180 226
342 226
342 209
356 209
1 2 14 0 0 4224 0 3 12 0 0 4
179 198
342 198
342 200
356 200
1 1 15 0 0 4224 0 4 12 0 0 4
178 171
342 171
342 191
356 191
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
