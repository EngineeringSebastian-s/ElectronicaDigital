CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files (x86)\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
13
13 Logic Switch~
5 136 293 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
45226.3 1
0
13 Logic Switch~
5 133 250 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
45226.3 0
0
13 Logic Switch~
5 134 216 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
45226.3 0
0
13 Logic Switch~
5 132 178 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
45226.3 0
0
5 4049~
219 699 292 0 2 22
0 7 8
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 2 0
1 U
8157 0 0
2
45226.3 0
0
5 4049~
219 697 260 0 2 22
0 6 9
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 2 0
1 U
5572 0 0
2
45226.3 0
0
5 4049~
219 698 229 0 2 22
0 5 10
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 2 0
1 U
8901 0 0
2
45226.3 0
0
5 4049~
219 732 206 0 2 22
0 4 11
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 2 0
1 U
7361 0 0
2
45226.3 0
0
5 4071~
219 865 243 0 3 22
0 13 8 12
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
4747 0 0
2
45226.3 0
0
5 4049~
219 732 164 0 2 22
0 2 14
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 2 0
1 U
972 0 0
2
45226.3 0
0
14 Logic Display~
6 905 165 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
45226.3 1
0
8 4-In OR~
219 809 225 0 5 22
0 14 11 10 9 13
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 1 0
1 U
9998 0 0
2
45226.3 0
0
6 74LS42
101 323 189 0 14 29
0 18 17 16 15 3 19 2 4 5
6 20 21 7 22
0
0 0 4848 0
6 74LS42
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
106 %D [%16bi %8bi %1i %2i %3i %4i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 11 10 9 7 6
5 4 3 2 1 12 13 14 15 11
10 9 7 6 5 4 3 2 1 0
65 0 0 512 0 0 0 0
1 U
3536 0 0
2
45226.3 0
0
18
7 1 2 0 0 4224 0 13 10 0 0 4
361 171
707 171
707 164
717 164
0 7 2 0 0 128 0 0 13 0 0 2
361 171
361 171
5 0 3 0 0 128 0 13 0 0 0 1
361 153
8 1 4 0 0 4240 0 13 8 0 0 4
361 180
705 180
705 206
717 206
9 1 5 0 0 4224 0 13 7 0 0 4
361 189
641 189
641 229
683 229
10 1 6 0 0 4224 0 13 6 0 0 4
361 198
606 198
606 260
682 260
13 1 7 0 0 8320 0 13 5 0 0 5
361 225
361 228
586 228
586 292
684 292
2 2 8 0 0 4224 0 5 9 0 0 3
720 292
852 292
852 252
2 4 9 0 0 4224 0 6 12 0 0 3
718 260
792 260
792 239
2 3 10 0 0 4224 0 7 12 0 0 4
719 229
793 229
793 230
792 230
2 2 11 0 0 8320 0 8 12 0 0 3
753 206
753 221
792 221
3 1 12 0 0 8320 0 9 11 0 0 3
898 243
905 243
905 183
1 5 13 0 0 8320 0 9 12 0 0 3
852 234
852 225
842 225
2 1 14 0 0 4224 0 10 12 0 0 4
753 164
793 164
793 212
792 212
1 4 15 0 0 4224 0 1 13 0 0 4
148 293
285 293
285 234
291 234
1 3 16 0 0 4224 0 2 13 0 0 4
145 250
263 250
263 225
291 225
1 2 17 0 0 4224 0 3 13 0 0 2
146 216
291 216
1 1 18 0 0 4224 0 4 13 0 0 4
144 178
283 178
283 207
291 207
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
