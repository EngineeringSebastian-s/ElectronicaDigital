CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
50 C:\Users\Edu\AppData\Local\Temp\IXP001.TMP\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
8
11 Multimeter~
205 659 273 0 17 21
0 3 10 11 5 0 0 0 0 0
78 79 32 68 65 84 65 32
0
0 0 16448 90
8 100.0Meg
-28 -19 28 -11
3 MM1
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
5130 0 0
2
5.90094e-315 0
0
8 Battery~
219 192 219 0 2 5
0 5 4
0
0 0 864 0
2 5V
15 -2 29 6
2 V1
16 -12 30 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
391 0 0
2
5.90094e-315 0
0
7 Ground~
168 562 622 0 1 3
0 12
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
3 GND
3124 0 0
2
5.90094e-315 0
0
8 2-In OR~
219 600 361 0 3 22
0 7 6 3
0
0 0 608 0
6 74LS32
-21 -24 21 -16
2 OR
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3421 0 0
2
5.90094e-315 0
0
9 2-In AND~
219 522 414 0 3 22
0 4 4 6
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 And
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
8157 0 0
2
5.90094e-315 0
0
9 2-In AND~
219 513 321 0 3 22
0 9 8 7
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 And
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
5572 0 0
2
5.90094e-315 0
0
9 Inverter~
13 387 380 0 2 22
0 4 8
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 notB
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
8901 0 0
2
5.90094e-315 0
0
9 Inverter~
13 385 337 0 2 22
0 4 9
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 notA
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
7361 0 0
2
5.90094e-315 0
0
17
0 0 0 0 0 16 0 0 0 0 0 2
239 444
239 444
0 0 0 0 0 0 0 0 0 0 0 2
321 442
321 442
0 0 0 0 0 4096 0 0 0 0 0 2
280 444
280 444
0 0 2 0 0 0 0 0 0 0 0 2
608 239
608 239
3 1 3 0 0 8320 0 4 1 0 0 4
633 361
683 361
683 304
676 304
0 0 4 0 0 4100 0 0 0 0 0 2
321 423
498 423
0 1 4 0 0 0 0 0 7 9 0 2
280 380
372 380
0 0 4 0 0 4 0 0 0 0 0 2
239 337
370 337
0 1 4 0 0 4096 0 0 5 11 0 3
280 239
280 405
498 405
0 1 4 0 0 16 0 0 8 11 0 3
239 239
239 337
370 337
2 2 4 0 0 0 0 2 5 0 0 5
192 230
192 239
321 239
321 423
498 423
1 4 5 0 0 8320 0 2 1 0 0 7
192 206
192 183
678 183
678 198
679 198
679 254
676 254
0 0 4 0 0 4228 0 0 0 0 0 2
280 405
498 405
3 2 6 0 0 8320 0 5 4 0 0 4
543 414
579 414
579 370
587 370
3 1 7 0 0 4224 0 6 4 0 0 4
534 321
579 321
579 352
587 352
2 2 8 0 0 4224 0 7 6 0 0 4
408 380
476 380
476 330
489 330
2 1 9 0 0 8320 0 8 6 0 0 5
406 337
406 296
481 296
481 312
489 312
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
227 211 254 232
236 217 244 232
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
267 212 292 233
275 218 283 233
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
306 208 333 229
315 215 323 230
1 C
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
