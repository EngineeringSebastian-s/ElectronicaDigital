CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
500 10 30 400 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files (x86)\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 607 41 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21104 0
2 5V
-6 -16 8 -8
6 toggle
-55 -5 -13 3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3472 0 0
2
45254.3 0
0
13 Logic Switch~
5 384 53 0 1 11
0 10
0
0 0 21232 0
2 0V
-6 -16 8 -8
3 set
-42 -7 -21 1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9998 0 0
2
45254.3 0
0
13 Logic Switch~
5 381 124 0 1 11
0 9
0
0 0 21232 0
2 0V
-6 -16 8 -8
5 reset
-49 -7 -14 1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3536 0 0
2
45254.3 0
0
13 Logic Switch~
5 382 82 0 1 11
0 13
0
0 0 21232 0
2 0V
-6 -16 8 -8
1 D
-20 -9 -13 -1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4597 0 0
2
45254.3 1
0
13 Logic Switch~
5 381 100 0 1 11
0 12
0
0 0 21104 0
2 0V
-6 -16 8 -8
3 clk
-34 -7 -13 1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3835 0 0
2
45254.3 0
0
13 Logic Switch~
5 380 177 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21104 0
2 5V
-6 -16 8 -8
3 clk
-34 -7 -13 1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3670 0 0
2
45254.3 0
0
13 Logic Switch~
5 381 159 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21232 0
2 5V
-6 -16 8 -8
1 D
-20 -9 -13 -1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5616 0 0
2
45254.3 0
0
2 +V
167 753 157 0 1 3
0 4
0
0 0 53488 270
3 10V
-11 -15 10 -7
2 V1
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9323 0 0
2
45254.3 0
0
2 +V
167 577 139 0 1 3
0 5
0
0 0 53488 90
3 10V
-11 -15 10 -7
2 V2
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
317 0 0
2
45254.3 0
0
14 Logic Display~
6 778 69 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3108 0 0
2
45254.3 0
0
14 NO PushButton~
191 665 148 0 2 5
0 7 2
0
0 0 4720 0
0
5 reset
-42 -9 -7 -1
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
4299 0 0
2
45254.3 1
0
7 Ground~
168 624 162 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9672 0 0
2
45254.3 0
0
7 Ground~
168 554 102 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7876 0 0
2
45254.3 0
0
14 NO PushButton~
191 589 88 0 2 5
0 6 2
0
0 0 4720 0
0
3 clk
-36 -9 -15 -1
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
6369 0 0
2
45254.3 0
0
6 JK RN~
219 691 104 0 6 22
0 3 6 3 7 17 8
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 2 0
1 U
9172 0 0
2
45254.3 0
0
14 Logic Display~
6 487 62 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7100 0 0
2
45254.3 0
0
5 4013~
219 417 118 0 6 22
0 10 13 12 9 18 11
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 1 0
1 U
3820 0 0
2
45254.3 0
0
12 D Flip-Flop~
219 415 195 0 4 9
0 15 14 19 16
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U2
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7678 0 0
2
45254.3 0
0
14 Logic Display~
6 487 141 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
961 0 0
2
45254.3 0
0
9 Resistor~
219 716 156 0 3 5
0 4 7 1
0
0 0 112 180
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3178 0 0
2
45254.3 0
0
9 Resistor~
219 657 294 0 2 5
0 20 21
0
0 0 112 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 512 0 0 0 0
1 R
3409 0 0
2
45254.3 0
0
9 Resistor~
219 623 119 0 3 5
0 5 6 1
0
0 0 112 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3951 0 0
2
45254.3 0
0
19
0 3 3 0 0 4096 0 0 15 6 0 3
652 87
652 105
667 105
1 1 4 0 0 4224 0 20 8 0 0 2
734 156
741 156
1 1 5 0 0 4224 0 22 9 0 0 2
623 137
588 137
0 2 6 0 0 4096 0 0 22 11 0 2
623 96
623 101
0 2 7 0 0 4224 0 0 20 8 0 2
690 156
698 156
1 1 3 0 0 8320 0 1 15 0 0 4
619 41
652 41
652 87
667 87
1 6 8 0 0 4224 0 10 15 0 0 2
778 87
715 87
1 4 7 0 0 8320 0 11 15 0 0 3
682 156
691 156
691 135
1 2 2 0 0 4224 0 12 11 0 0 2
624 156
648 156
1 2 2 0 0 128 0 13 14 0 0 2
554 96
572 96
1 2 6 0 0 4224 0 14 15 0 0 2
606 96
660 96
1 4 9 0 0 4224 0 3 17 0 0 2
393 124
417 124
1 1 10 0 0 8320 0 17 2 0 0 4
417 61
417 54
396 54
396 53
1 6 11 0 0 8320 0 16 17 0 0 3
487 80
487 82
441 82
1 3 12 0 0 0 0 5 17 0 0 2
393 100
393 100
1 2 13 0 0 4224 0 4 17 0 0 2
394 82
393 82
1 2 14 0 0 4224 0 6 18 0 0 2
392 177
391 177
1 1 15 0 0 4224 0 7 18 0 0 2
393 159
391 159
1 4 16 0 0 4224 0 19 18 0 0 2
487 159
439 159
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
