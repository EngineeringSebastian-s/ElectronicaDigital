CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 90 30 200 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files (x86)\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
41
13 Logic Switch~
5 127 828 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-28 -3 -14 5
2 S2
-28 -13 -14 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90099e-315 0
0
13 Logic Switch~
5 71 520 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
6 Select
-20 -26 22 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.90099e-315 0
0
13 Logic Switch~
5 74 687 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.90099e-315 5.32571e-315
0
13 Logic Switch~
5 74 718 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.90099e-315 5.30499e-315
0
13 Logic Switch~
5 75 754 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
5.90099e-315 5.26354e-315
0
13 Logic Switch~
5 76 788 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.90099e-315 0
0
13 Logic Switch~
5 73 658 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
5.90099e-315 0
0
13 Logic Switch~
5 72 624 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
5.90099e-315 0
0
13 Logic Switch~
5 71 589 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4747 0 0
2
5.90099e-315 0
0
13 Logic Switch~
5 71 557 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
972 0 0
2
5.90099e-315 0
0
13 Logic Switch~
5 121 326 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-32 -3 -18 5
2 A2
-29 -15 -15 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
5.90099e-315 5.3568e-315
0
13 Logic Switch~
5 122 385 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-32 -3 -18 5
2 A0
-29 -15 -15 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
5.90099e-315 5.34643e-315
0
13 Logic Switch~
5 121 354 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-30 -1 -16 7
2 A1
-30 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
5.90099e-315 5.32571e-315
0
13 Logic Switch~
5 124 441 0 1 11
0 22
0
0 0 21360 0
2 0V
-32 -3 -18 5
2 S0
-29 -15 -15 -7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4597 0 0
2
5.90099e-315 5.30499e-315
0
13 Logic Switch~
5 123 410 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-30 -1 -16 7
2 S1
-30 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3835 0 0
2
5.90099e-315 5.26354e-315
0
13 Logic Switch~
5 120 295 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-30 -1 -16 7
2 A3
-30 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3670 0 0
2
5.90099e-315 0
0
13 Logic Switch~
5 154 246 0 1 11
0 37
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5616 0 0
2
5.90099e-315 0
0
13 Logic Switch~
5 153 209 0 10 11
0 36 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9323 0 0
2
5.90099e-315 0
0
13 Logic Switch~
5 153 175 0 1 11
0 39
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 S
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
317 0 0
2
5.90099e-315 0
0
14 Logic Display~
6 414 863 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
5.90099e-315 0
0
5 4071~
219 369 884 0 3 22
0 5 4 3
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
4299 0 0
2
5.90099e-315 0
0
5 4049~
219 319 825 0 2 22
0 6 7
0
0 0 624 270
4 4049
-7 -24 21 -16
3 U3F
-22 -24 -1 -16
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 3 0
1 U
9672 0 0
2
5.90099e-315 0
0
7 74LS153
119 279 882 0 14 29
0 43 44 45 46 47 48 49 50 51
52 7 6 5 4
0
0 0 4848 0
6 74F153
-21 -60 21 -52
2 U8
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 512 1 0 0 0
1 U
7876 0 0
2
5.90099e-315 0
0
7 Ground~
168 248 721 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6369 0 0
2
5.90099e-315 0
0
7 74LS157
122 285 622 0 14 29
0 16 13 9 12 8 11 14 10 15
2 20 19 18 17
0
0 0 4848 0
6 74F157
-21 -60 21 -52
2 U7
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
9172 0 0
2
5.90099e-315 5.26354e-315
0
12 Hex Display~
7 405 557 0 18 19
10 17 18 19 20 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
7100 0 0
2
5.90099e-315 0
0
14 Logic Display~
6 475 351 0 1 2
10 27
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
5.90099e-315 0
0
5 4049~
219 262 405 0 2 22
0 22 28
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3E
2 -13 23 -5
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
7678 0 0
2
5.90099e-315 0
0
5 4049~
219 255 341 0 2 22
0 23 29
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3D
3 -16 24 -8
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
961 0 0
2
5.90099e-315 0
0
5 4049~
219 254 311 0 2 22
0 22 30
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3C
3 -16 24 -8
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
3178 0 0
2
5.90099e-315 0
0
5 4049~
219 254 285 0 2 22
0 23 31
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
2 -17 23 -9
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
3409 0 0
2
5.90099e-315 0
0
8 4-In OR~
219 422 381 0 5 22
0 35 34 33 32 27
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
3951 0 0
2
5.90099e-315 0
0
5 7415~
219 318 458 0 4 22
0 23 22 21 32
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 5 0
1 U
8885 0 0
2
5.90099e-315 0
0
5 7415~
219 316 410 0 4 22
0 23 28 24 33
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 4 0
1 U
3780 0 0
2
5.90099e-315 0
0
5 7415~
219 315 357 0 4 22
0 29 22 25 34
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 4 0
1 U
9265 0 0
2
5.90099e-315 0
0
5 7415~
219 313 308 0 4 22
0 31 30 26 35
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 4 0
1 U
9442 0 0
2
5.90099e-315 0
0
14 Logic Display~
6 462 186 0 1 2
10 38
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
5.90099e-315 0
0
5 4049~
219 250 173 0 2 22
0 39 40
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
9968 0 0
2
5.90099e-315 0
0
5 4071~
219 374 213 0 3 22
0 42 41 38
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
9281 0 0
2
5.90099e-315 0
0
5 4081~
219 314 239 0 3 22
0 39 36 41
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
8464 0 0
2
5.90099e-315 0
0
5 4081~
219 314 182 0 3 22
0 40 37 42
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
7168 0 0
2
5.90099e-315 0
0
49
1 3 3 0 0 8320 0 20 21 0 0 3
414 881
414 884
402 884
2 14 4 0 0 8320 0 21 23 0 0 3
356 893
356 909
311 909
1 13 5 0 0 8320 0 21 23 0 0 3
356 875
356 864
311 864
0 12 6 0 0 12416 0 0 23 5 0 5
322 799
322 798
337 798
337 927
317 927
1 1 6 0 0 0 0 1 22 0 0 5
139 828
243 828
243 799
322 799
322 807
2 11 7 0 0 8320 0 22 23 0 0 3
322 843
322 846
317 846
1 5 8 0 0 4224 0 4 25 0 0 4
86 718
215 718
215 622
253 622
1 3 9 0 0 4224 0 3 25 0 0 4
86 687
205 687
205 604
253 604
1 8 10 0 0 4224 0 7 25 0 0 4
85 658
230 658
230 649
253 649
1 6 11 0 0 8320 0 8 25 0 0 5
84 624
84 630
239 630
239 631
253 631
1 4 12 0 0 4224 0 9 25 0 0 4
83 589
234 589
234 613
253 613
1 2 13 0 0 4224 0 10 25 0 0 4
83 557
239 557
239 595
253 595
1 7 14 0 0 4224 0 5 25 0 0 4
87 754
223 754
223 640
253 640
1 9 15 0 0 4224 0 6 25 0 0 4
88 788
234 788
234 658
253 658
1 1 16 0 0 4224 0 2 25 0 0 4
83 520
246 520
246 586
253 586
1 10 2 0 0 8320 0 24 25 0 0 5
248 715
246 715
246 666
247 666
247 667
14 1 17 0 0 4224 0 25 26 0 0 3
317 658
414 658
414 581
13 2 18 0 0 4224 0 25 26 0 0 3
317 640
408 640
408 581
12 3 19 0 0 4224 0 25 26 0 0 3
317 622
402 622
402 581
11 4 20 0 0 4224 0 25 26 0 0 3
317 604
396 604
396 581
1 3 21 0 0 8320 0 16 33 0 0 4
132 295
144 295
144 467
294 467
0 2 22 0 0 12288 0 0 33 31 0 4
199 441
226 441
226 458
294 458
0 1 23 0 0 8192 0 0 33 32 0 3
231 410
231 449
294 449
1 3 24 0 0 12416 0 11 34 0 0 4
133 326
152 326
152 419
292 419
0 1 22 0 0 0 0 0 28 31 0 3
199 401
247 401
247 405
0 1 23 0 0 0 0 0 34 32 0 4
231 391
288 391
288 401
292 401
1 3 25 0 0 8320 0 13 35 0 0 3
133 354
133 366
291 366
0 2 22 0 0 4096 0 0 35 31 0 2
199 357
291 357
0 1 23 0 0 0 0 0 29 32 0 2
231 341
240 341
1 3 26 0 0 12416 0 12 36 0 0 5
134 385
158 385
158 326
289 326
289 317
1 1 22 0 0 8320 0 14 30 0 0 4
136 441
199 441
199 311
239 311
1 1 23 0 0 8320 0 15 31 0 0 4
135 410
231 410
231 285
239 285
1 5 27 0 0 8320 0 27 32 0 0 4
475 369
475 380
455 380
455 381
2 2 28 0 0 8320 0 28 34 0 0 3
283 405
283 410
292 410
2 1 29 0 0 8320 0 29 35 0 0 3
276 341
276 348
291 348
2 2 30 0 0 4224 0 30 36 0 0 3
275 311
289 311
289 308
2 1 31 0 0 4224 0 31 36 0 0 3
275 285
289 285
289 299
4 4 32 0 0 8320 0 33 32 0 0 4
339 458
392 458
392 395
405 395
4 3 33 0 0 4224 0 34 32 0 0 4
337 410
386 410
386 386
405 386
4 2 34 0 0 4224 0 35 32 0 0 4
336 357
392 357
392 377
405 377
4 1 35 0 0 4224 0 36 32 0 0 4
334 308
397 308
397 368
405 368
1 2 36 0 0 12416 0 18 40 0 0 4
165 209
175 209
175 248
290 248
1 2 37 0 0 16512 0 17 41 0 0 5
166 246
166 221
200 221
200 191
290 191
1 3 38 0 0 8320 0 37 39 0 0 3
462 204
462 213
407 213
0 1 39 0 0 8320 0 0 40 46 0 3
206 173
206 230
290 230
1 1 39 0 0 0 0 19 38 0 0 3
165 175
165 173
235 173
2 1 40 0 0 4224 0 38 41 0 0 2
271 173
290 173
2 3 41 0 0 4224 0 39 40 0 0 4
361 222
338 222
338 239
335 239
1 3 42 0 0 4224 0 39 41 0 0 3
361 204
335 204
335 182
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
