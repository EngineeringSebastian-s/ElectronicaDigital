CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 40 30 120 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
47
13 Logic Switch~
5 48 83 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21088 0
2 5V
-6 -16 8 -8
2 S1
-13 -17 1 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7376 0 0
2
5.90101e-315 5.47595e-315
0
13 Logic Switch~
5 64 297 0 1 11
0 17
0
0 0 21088 0
2 0V
-6 -16 8 -8
2 B3
-27 -4 -13 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9156 0 0
2
5.90101e-315 5.47207e-315
0
13 Logic Switch~
5 60 191 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21088 0
2 5V
-6 -16 8 -8
2 A3
-26 -4 -12 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5776 0 0
2
5.90101e-315 5.47077e-315
0
13 Logic Switch~
5 48 112 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21088 0
2 5V
-6 -16 8 -8
2 S0
-13 -17 1 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7207 0 0
2
5.90101e-315 5.46818e-315
0
13 Logic Switch~
5 60 233 0 1 11
0 14
0
0 0 21088 0
2 0V
-6 -16 8 -8
2 A1
-27 -4 -13 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4459 0 0
2
5.90101e-315 5.46559e-315
0
13 Logic Switch~
5 60 214 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21088 0
2 5V
-6 -16 8 -8
2 A2
-26 -4 -12 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3760 0 0
2
5.90101e-315 5.463e-315
0
13 Logic Switch~
5 61 252 0 1 11
0 12
0
0 0 21088 0
2 0V
-6 -16 8 -8
2 A0
-27 -4 -13 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
754 0 0
2
5.90101e-315 5.46041e-315
0
13 Logic Switch~
5 65 317 0 1 11
0 15
0
0 0 21088 0
2 0V
-6 -16 8 -8
2 B2
-27 -4 -13 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9767 0 0
2
5.90101e-315 5.45782e-315
0
13 Logic Switch~
5 66 337 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21088 0
2 5V
-6 -16 8 -8
2 B1
-27 -4 -13 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7978 0 0
2
5.90101e-315 5.45523e-315
0
13 Logic Switch~
5 67 362 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21088 0
2 5V
-6 -16 8 -8
2 B0
-27 -4 -13 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3142 0 0
2
5.90101e-315 5.45264e-315
0
5 4071~
219 217 757 0 3 22
0 12 11 19
0
0 0 96 0
4 4071
-7 -24 21 -16
4 U14D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 6 0
1 U
3284 0 0
2
5.90101e-315 0
0
5 4071~
219 216 719 0 3 22
0 14 13 20
0
0 0 96 0
4 4071
-7 -24 21 -16
4 U14C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 6 0
1 U
659 0 0
2
5.90101e-315 0
0
5 4071~
219 214 682 0 3 22
0 16 15 21
0
0 0 96 0
4 4071
-7 -24 21 -16
4 U14B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
3800 0 0
2
5.90101e-315 0
0
5 4071~
219 213 643 0 3 22
0 18 17 22
0
0 0 96 0
4 4071
-7 -24 21 -16
4 U14A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
6792 0 0
2
5.90101e-315 0
0
7 Ground~
168 633 589 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3701 0 0
2
5.90101e-315 0
0
5 4081~
219 213 591 0 3 22
0 12 11 27
0
0 0 96 0
4 4081
-7 -24 21 -16
4 U13D
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
6316 0 0
2
5.90101e-315 0
0
5 4081~
219 212 556 0 3 22
0 14 13 28
0
0 0 96 0
4 4081
-7 -24 21 -16
4 U13C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
8734 0 0
2
5.90101e-315 0
0
5 4081~
219 212 518 0 3 22
0 16 15 29
0
0 0 96 0
4 4081
-7 -24 21 -16
4 U13B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
7988 0 0
2
5.90101e-315 0
0
5 4081~
219 211 483 0 3 22
0 18 17 30
0
0 0 96 0
4 4081
-7 -24 21 -16
4 U13A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
3217 0 0
2
5.90101e-315 0
0
7 74LS157
122 673 539 0 14 29
0 31 22 30 21 29 20 28 19 27
2 26 25 24 23
0
0 0 4832 0
6 74F157
-21 -60 21 -52
3 U12
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3965 0 0
2
5.90101e-315 0
0
7 Ground~
168 861 469 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8239 0 0
2
5.90101e-315 5.47466e-315
0
7 74LS157
122 900 416 0 14 29
0 10 26 35 25 34 24 33 23 32
2 39 38 37 36
0
0 0 4832 0
6 74F157
-21 -60 21 -52
3 U11
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
828 0 0
2
5.90101e-315 5.47336e-315
0
2 +V
167 626 348 0 1 3
0 41
0
0 0 53472 90
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6187 0 0
2
5.90101e-315 5.45005e-315
0
9 CC 7-Seg~
183 1070 163 0 18 19
10 9 8 7 6 5 4 3 124 125
1 0 0 0 1 1 1 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7107 0 0
2
5.90101e-315 5.44746e-315
0
7 Ground~
168 749 347 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6433 0 0
2
5.90101e-315 5.44228e-315
0
7 74LS157
122 790 287 0 14 29
0 49 48 44 47 43 46 42 45 40
2 35 34 33 32
0
0 0 4832 0
6 74F157
-21 -60 21 -52
2 U9
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
8559 0 0
2
5.90101e-315 5.43969e-315
0
9 Inverter~
13 569 315 0 2 22
0 40 50
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U8A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3674 0 0
2
5.90101e-315 5.4371e-315
0
9 Inverter~
13 583 273 0 2 22
0 43 52
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U3F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
5697 0 0
2
5.90101e-315 5.43451e-315
0
9 Inverter~
13 569 290 0 2 22
0 42 51
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U3E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
3805 0 0
2
5.90101e-315 5.43192e-315
0
9 Inverter~
13 578 250 0 2 22
0 44 53
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
5219 0 0
2
5.90101e-315 5.42933e-315
0
7 Ground~
168 621 323 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3795 0 0
2
5.90101e-315 5.42414e-315
0
6 74LS83
105 670 302 0 14 29
0 53 52 51 50 2 2 2 2 41
48 47 46 45 126
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U7
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3637 0 0
2
5.90101e-315 5.41896e-315
0
9 CC 7-Seg~
183 1004 163 0 18 19
10 127 128 129 130 131 132 49 133 10
2 2 2 2 2 2 1 2 1
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP2
-72 -17 -37 -9
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3226 0 0
2
5.90101e-315 5.41378e-315
0
9 2-In AND~
219 489 150 0 3 22
0 31 44 49
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6966 0 0
2
5.90101e-315 5.4086e-315
0
12 Hex Display~
7 226 153 0 18 19
10 11 13 15 17 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
1 B
-4 -38 3 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9796 0 0
2
5.90101e-315 5.40342e-315
0
12 Hex Display~
7 187 154 0 18 19
10 12 14 16 18 0 0 0 0 0
0 1 0 0 1 1 1 0 12
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
1 A
-4 -38 3 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5952 0 0
2
5.90101e-315 5.39824e-315
0
9 Inverter~
13 208 278 0 2 22
0 17 54
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
3649 0 0
2
5.90101e-315 5.39306e-315
0
2 +V
167 206 378 0 1 3
0 63
0
0 0 53472 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3716 0 0
2
5.90101e-315 5.38788e-315
0
7 Ground~
168 224 370 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4797 0 0
2
5.90101e-315 5.37752e-315
0
9 Inverter~
13 206 324 0 2 22
0 13 65
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
4681 0 0
2
5.90101e-315 5.36716e-315
0
9 Inverter~
13 206 299 0 2 22
0 15 66
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U2F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
9730 0 0
2
5.90101e-315 5.3568e-315
0
9 Inverter~
13 206 348 0 2 22
0 11 64
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
9874 0 0
2
5.90101e-315 5.34643e-315
0
6 74LS83
105 283 335 0 14 29
0 54 66 65 64 2 2 2 2 63
56 57 58 55 134
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
364 0 0
2
5.90101e-315 5.32571e-315
0
7 74LS157
122 384 329 0 14 29
0 31 56 17 57 15 58 13 55 11
2 59 60 61 62
0
0 0 4832 0
6 74F157
-21 -60 21 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3656 0 0
2
5.90101e-315 5.30499e-315
0
7 Ground~
168 451 373 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3131 0 0
2
5.90101e-315 5.26354e-315
0
6 74LS83
105 477 271 0 14 29
0 18 16 14 12 59 60 61 62 2
44 43 42 40 135
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
6772 0 0
2
5.90101e-315 0
0
12 DEC_BCH_7SEG
94 1000 431 0 11 23
0 39 38 37 36 3 4 5 6 7
8 9
12 DEC_BCH_7SEG
1 0 4736 0
0
3 U15
-11 -55 10 -47
0
0
0
0
0
0
23

0 1 2 3 4 10 11 12 13 14
15 16 1 2 3 4 10 11 12 13
14 15 16 0
0 0 0 0 1 0 0 0
1 U
9557 0 0
2
5.90097e-315 0
0
115
5 7 3 0 0 8320 0 47 24 0 0 3
1033 458
1085 458
1085 199
6 6 4 0 0 8320 0 47 24 0 0 3
1033 449
1079 449
1079 199
7 5 5 0 0 8320 0 47 24 0 0 3
1033 440
1073 440
1073 199
8 4 6 0 0 8320 0 47 24 0 0 3
1033 431
1067 431
1067 199
9 3 7 0 0 8320 0 47 24 0 0 3
1033 422
1061 422
1061 199
10 2 8 0 0 8320 0 47 24 0 0 3
1033 413
1055 413
1055 199
11 1 9 0 0 8320 0 47 24 0 0 3
1033 404
1049 404
1049 199
0 9 10 0 0 4096 0 0 33 42 0 3
863 100
1004 100
1004 121
0 2 11 0 0 4096 0 0 11 21 0 3
115 600
115 766
204 766
0 1 12 0 0 4096 0 0 11 22 0 3
122 582
122 748
204 748
0 2 13 0 0 4096 0 0 12 23 0 3
131 565
131 728
203 728
0 1 14 0 0 4096 0 0 12 24 0 3
138 547
138 710
203 710
0 2 15 0 0 4096 0 0 13 25 0 3
148 527
148 691
201 691
0 1 16 0 0 4096 0 0 13 26 0 3
154 509
154 673
201 673
0 2 17 0 0 4096 0 0 14 27 0 3
168 492
168 652
200 652
0 1 18 0 0 4096 0 0 14 28 0 3
178 474
178 634
200 634
3 8 19 0 0 4224 0 11 20 0 0 4
250 757
609 757
609 566
641 566
3 6 20 0 0 4224 0 12 20 0 0 4
249 719
602 719
602 548
641 548
3 4 21 0 0 4224 0 13 20 0 0 4
247 682
592 682
592 530
641 530
3 2 22 0 0 4224 0 14 20 0 0 4
246 643
586 643
586 512
641 512
0 2 11 0 0 4224 0 0 16 106 0 3
85 362
85 600
189 600
0 1 12 0 0 4224 0 0 16 115 0 3
78 252
78 582
189 582
0 2 13 0 0 4224 0 0 17 107 0 3
92 337
92 565
188 565
0 1 14 0 0 4096 0 0 17 114 0 3
100 224
100 547
188 547
0 2 15 0 0 4224 0 0 18 90 0 3
108 317
108 527
188 527
0 1 16 0 0 4224 0 0 18 113 0 3
113 203
113 509
188 509
0 2 17 0 0 4224 0 0 19 84 0 3
125 297
125 492
187 492
0 1 18 0 0 4224 0 0 19 87 0 3
133 191
133 474
187 474
14 8 23 0 0 8320 0 20 22 0 0 4
705 575
825 575
825 443
868 443
13 6 24 0 0 8320 0 20 22 0 0 4
705 557
835 557
835 425
868 425
0 13 24 0 0 0 0 0 20 0 0 3
694 558
694 557
705 557
12 4 25 0 0 8320 0 20 22 0 0 4
705 539
816 539
816 407
868 407
11 2 26 0 0 8320 0 20 22 0 0 4
705 521
806 521
806 389
868 389
1 10 2 0 0 8192 0 15 20 0 0 3
633 583
633 584
635 584
3 9 27 0 0 4224 0 16 20 0 0 4
234 591
627 591
627 575
641 575
3 7 28 0 0 4224 0 17 20 0 0 4
233 556
627 556
627 557
641 557
3 5 29 0 0 4224 0 18 20 0 0 4
233 518
622 518
622 539
641 539
3 3 30 0 0 4224 0 19 20 0 0 4
232 483
627 483
627 521
641 521
0 1 31 0 0 8320 0 0 20 88 0 4
143 112
143 450
641 450
641 503
1 0 12 0 0 0 0 36 0 0 115 4
196 178
196 228
197 228
197 233
0 1 31 0 0 0 0 0 34 88 0 2
332 141
465 141
1 1 10 0 0 8320 0 1 22 0 0 5
60 83
60 81
863 81
863 380
868 380
1 10 2 0 0 0 0 21 22 0 0 3
861 463
861 461
862 461
14 9 32 0 0 8320 0 26 22 0 0 4
822 323
839 323
839 452
868 452
13 7 33 0 0 8320 0 26 22 0 0 4
822 305
844 305
844 434
868 434
12 5 34 0 0 8320 0 26 22 0 0 4
822 287
849 287
849 416
868 416
11 3 35 0 0 8320 0 26 22 0 0 4
822 269
854 269
854 398
868 398
14 4 36 0 0 4224 0 22 47 0 0 4
932 452
963 452
963 431
967 431
13 3 37 0 0 4224 0 22 47 0 0 4
932 434
960 434
960 422
967 422
12 2 38 0 0 4224 0 22 47 0 0 4
932 416
960 416
960 413
967 413
11 1 39 0 0 4224 0 22 47 0 0 4
932 398
960 398
960 404
967 404
0 9 40 0 0 8320 0 0 26 72 0 5
519 315
519 414
738 414
738 323
758 323
1 0 2 0 0 8192 0 31 0 0 55 3
621 317
621 316
638 316
7 8 2 0 0 0 0 32 32 0 0 2
638 320
638 329
6 7 2 0 0 0 0 32 32 0 0 2
638 311
638 320
5 6 2 0 0 0 0 32 32 0 0 2
638 302
638 311
1 9 41 0 0 4224 0 23 32 0 0 3
637 346
637 347
638 347
10 1 2 0 0 0 0 26 25 0 0 3
752 332
749 332
749 341
7 0 42 0 0 12416 0 26 0 0 73 5
758 305
732 305
732 405
527 405
527 280
0 5 43 0 0 8320 0 0 26 74 0 5
543 271
543 393
727 393
727 287
758 287
0 3 44 0 0 8320 0 0 26 75 0 5
535 250
535 377
719 377
719 269
758 269
13 8 45 0 0 12416 0 32 26 0 0 5
702 320
705 320
705 317
758 317
758 314
12 6 46 0 0 16512 0 32 26 0 0 5
702 311
702 312
713 312
713 296
758 296
11 4 47 0 0 12416 0 32 26 0 0 4
702 302
710 302
710 278
758 278
10 2 48 0 0 12416 0 32 26 0 0 4
702 293
705 293
705 260
758 260
0 1 49 0 0 4096 0 0 26 76 0 3
743 219
743 251
758 251
2 0 44 0 0 0 0 34 0 0 75 5
465 159
460 159
460 189
535 189
535 250
2 4 50 0 0 12416 0 27 32 0 0 4
590 315
604 315
604 293
638 293
2 3 51 0 0 12416 0 29 32 0 0 4
590 290
598 290
598 284
638 284
2 2 52 0 0 12416 0 28 32 0 0 4
604 273
607 273
607 275
638 275
2 1 53 0 0 4224 0 30 32 0 0 4
599 250
620 250
620 266
638 266
13 1 40 0 0 0 0 46 27 0 0 4
509 289
514 289
514 315
554 315
12 1 42 0 0 0 0 46 29 0 0 3
509 280
554 280
554 290
11 1 43 0 0 0 0 46 28 0 0 3
509 271
568 271
568 273
10 1 44 0 0 0 0 46 30 0 0 4
509 262
516 262
516 250
563 250
3 7 49 0 0 12416 0 34 33 0 0 5
510 150
587 150
587 219
1019 219
1019 199
4 0 17 0 0 0 0 35 0 0 85 5
217 177
217 243
162 243
162 264
152 264
3 0 15 0 0 0 0 35 0 0 108 4
223 177
223 247
177 247
177 289
2 0 13 0 0 0 0 35 0 0 107 4
229 177
229 254
182 254
182 324
1 1 11 0 0 0 0 35 42 0 0 5
235 177
235 258
187 258
187 348
191 348
2 0 14 0 0 0 0 36 0 0 114 2
190 178
190 224
3 0 16 0 0 0 0 36 0 0 113 2
184 178
184 201
4 0 18 0 0 0 0 36 0 0 87 2
178 178
178 185
3 1 17 0 0 0 0 44 2 0 0 6
352 311
326 311
326 442
152 442
152 297
76 297
1 1 17 0 0 0 0 2 37 0 0 6
76 297
152 297
152 264
162 264
162 278
193 278
2 1 54 0 0 8320 0 37 43 0 0 4
229 278
231 278
231 299
251 299
1 1 18 0 0 0 0 3 46 0 0 6
72 191
178 191
178 185
431 185
431 235
445 235
1 1 31 0 0 0 0 4 44 0 0 4
60 112
332 112
332 293
352 293
10 0 2 0 0 8320 0 44 0 0 112 5
346 374
346 418
434 418
434 341
443 341
1 5 15 0 0 0 0 8 44 0 0 6
77 317
159 317
159 432
332 432
332 329
352 329
0 7 13 0 0 0 0 0 44 107 0 5
175 324
175 425
337 425
337 347
352 347
1 9 11 0 0 0 0 42 44 0 0 6
191 348
187 348
187 413
342 413
342 365
352 365
13 8 55 0 0 12416 0 43 44 0 0 4
315 353
321 353
321 356
352 356
2 10 56 0 0 4224 0 44 43 0 0 4
352 302
318 302
318 326
315 326
4 11 57 0 0 4224 0 44 43 0 0 4
352 320
322 320
322 335
315 335
12 6 58 0 0 12416 0 43 44 0 0 4
315 344
322 344
322 338
352 338
11 5 59 0 0 8320 0 44 46 0 0 4
416 311
417 311
417 271
445 271
12 6 60 0 0 8320 0 44 46 0 0 4
416 329
422 329
422 280
445 280
13 7 61 0 0 8320 0 44 46 0 0 4
416 347
427 347
427 289
445 289
14 8 62 0 0 8320 0 44 46 0 0 4
416 365
430 365
430 298
445 298
9 1 63 0 0 12416 0 43 38 0 0 4
251 380
237 380
237 387
206 387
8 0 2 0 0 0 0 43 0 0 105 2
251 362
238 362
7 0 2 0 0 0 0 43 0 0 105 2
251 353
238 353
6 0 2 0 0 0 0 43 0 0 105 2
251 344
238 344
5 1 2 0 0 0 0 43 39 0 0 4
251 335
238 335
238 364
224 364
1 1 11 0 0 0 0 42 10 0 0 4
191 348
181 348
181 362
79 362
1 1 13 0 0 0 0 40 9 0 0 4
191 324
168 324
168 337
78 337
1 1 15 0 0 0 0 41 8 0 0 5
191 299
191 289
159 289
159 317
77 317
4 2 64 0 0 4224 0 43 42 0 0 4
251 326
229 326
229 348
227 348
3 2 65 0 0 4224 0 43 40 0 0 4
251 317
225 317
225 324
227 324
2 2 66 0 0 4224 0 43 41 0 0 4
251 308
225 308
225 299
227 299
1 9 2 0 0 0 0 45 46 0 0 5
451 367
451 341
443 341
443 316
445 316
1 2 16 0 0 0 0 6 46 0 0 7
72 214
72 203
184 203
184 201
419 201
419 244
445 244
1 3 14 0 0 8320 0 5 46 0 0 5
72 233
72 224
413 224
413 253
445 253
1 4 12 0 0 0 0 7 46 0 0 6
73 252
148 252
148 233
406 233
406 262
445 262
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
