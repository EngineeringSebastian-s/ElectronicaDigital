CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
30 20 30 200 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
50 C:\Users\Edu\AppData\Local\Temp\IXP001.TMP\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
24
13 Logic Switch~
5 216 61 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9172 0 0
2
45219.3 1
0
13 Logic Switch~
5 213 103 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7100 0 0
2
45219.3 3
0
13 Logic Switch~
5 212 143 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3820 0 0
2
45219.3 2
0
13 Logic Switch~
5 211 176 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7678 0 0
2
45219.3 1
0
13 Logic Switch~
5 211 209 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
961 0 0
2
45219.3 0
0
13 Logic Switch~
5 208 356 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3178 0 0
2
45219.3 0
0
13 Logic Switch~
5 208 323 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3409 0 0
2
45219.3 0
0
13 Logic Switch~
5 209 290 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3951 0 0
2
45219.3 0
0
13 Logic Switch~
5 210 250 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8885 0 0
2
45219.3 0
0
5 4069~
219 284 66 0 2 22
0 3 2
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U4A
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
3780 0 0
2
45219.3 0
0
5 4069~
219 279 210 0 2 22
0 8 7
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U3F
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 6 2 0
1 U
9265 0 0
2
45219.3 7
0
5 4069~
219 281 108 0 2 22
0 11 4
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U3E
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 5 2 0
1 U
9442 0 0
2
45219.3 6
0
5 4069~
219 280 141 0 2 22
0 10 5
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U3D
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 4 2 0
1 U
9424 0 0
2
45219.3 5
0
5 4069~
219 280 177 0 2 22
0 9 6
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U3C
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 3 2 0
1 U
9968 0 0
2
45219.3 4
0
5 4069~
219 277 324 0 2 22
0 17 14
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 2 2 0
1 U
9281 0 0
2
45219.3 3
0
5 4069~
219 277 288 0 2 22
0 18 13
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 1 2 0
1 U
8464 0 0
2
45219.3 2
0
5 4069~
219 278 255 0 2 22
0 19 12
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U2F
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 6 1 0
1 U
7168 0 0
2
45219.3 1
0
5 4069~
219 276 357 0 2 22
0 16 15
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U2E
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 5 1 0
1 U
3171 0 0
2
45219.3 0
0
12 Hex Display~
7 639 262 0 16 19
10 24 25 26 27 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
4139 0 0
2
45219.3 0
0
5 4069~
219 477 256 0 2 22
0 23 27
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U2A
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
6435 0 0
2
45219.3 3
0
5 4069~
219 476 289 0 2 22
0 22 26
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U2B
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 2 1 0
1 U
5283 0 0
2
45219.3 2
0
5 4069~
219 476 325 0 2 22
0 21 25
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U2C
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 3 1 0
1 U
6874 0 0
2
45219.3 1
0
5 4069~
219 475 358 0 2 22
0 20 24
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U2D
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 4 1 0
1 U
5305 0 0
2
45219.3 0
0
5 74147
219 379 306 0 13 27
0 2 4 5 6 7 12 13 14 15
20 21 22 23
0
0 0 4848 0
5 74147
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
121 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
27

0 10 5 4 3 2 1 13 12 11
9 7 6 14 10 5 4 3 2 1
13 12 11 9 7 6 14 0
65 0 0 0 0 0 0 0
1 U
34 0 0
2
45219.3 0
0
26
2 1 2 0 0 8320 0 10 24 0 0 4
305 66
346 66
346 270
341 270
1 1 3 0 0 4224 0 1 10 0 0 4
228 61
261 61
261 66
269 66
2 2 4 0 0 8320 0 12 24 0 0 4
302 108
339 108
339 279
341 279
2 3 5 0 0 8336 0 13 24 0 0 4
301 141
334 141
334 288
341 288
2 4 6 0 0 8320 0 14 24 0 0 4
301 177
330 177
330 297
341 297
2 5 7 0 0 12416 0 11 24 0 0 5
300 210
300 209
324 209
324 306
341 306
1 1 8 0 0 4224 0 5 11 0 0 4
223 209
256 209
256 210
264 210
1 1 9 0 0 4224 0 4 14 0 0 4
223 176
257 176
257 177
265 177
1 1 10 0 0 4224 0 3 13 0 0 4
224 143
257 143
257 141
265 141
1 1 11 0 0 4224 0 2 12 0 0 4
225 103
258 103
258 108
266 108
2 6 12 0 0 8320 0 17 24 0 0 4
299 255
319 255
319 315
341 315
2 7 13 0 0 8320 0 16 24 0 0 4
298 288
314 288
314 324
341 324
2 8 14 0 0 8320 0 15 24 0 0 5
298 324
298 331
333 331
333 333
341 333
2 9 15 0 0 4224 0 18 24 0 0 4
297 357
333 357
333 342
341 342
1 1 16 0 0 4224 0 6 18 0 0 4
220 356
253 356
253 357
261 357
1 1 17 0 0 4224 0 7 15 0 0 4
220 323
254 323
254 324
262 324
1 1 18 0 0 4224 0 8 16 0 0 4
221 290
254 290
254 288
262 288
1 1 19 0 0 4224 0 9 17 0 0 4
222 250
255 250
255 255
263 255
10 1 20 0 0 8320 0 24 23 0 0 4
417 315
447 315
447 358
460 358
11 1 21 0 0 4224 0 24 22 0 0 4
417 306
453 306
453 325
461 325
12 1 22 0 0 4224 0 24 21 0 0 5
417 297
453 297
453 292
461 292
461 289
13 1 23 0 0 4224 0 24 20 0 0 4
417 288
454 288
454 256
462 256
2 1 24 0 0 4224 0 23 19 0 0 3
496 358
648 358
648 286
2 2 25 0 0 4224 0 22 19 0 0 3
497 325
642 325
642 286
2 3 26 0 0 4224 0 21 19 0 0 5
497 289
604 289
604 301
636 301
636 286
2 4 27 0 0 4224 0 20 19 0 0 5
498 256
609 256
609 296
630 296
630 286
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
