CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
10 60 30 200 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
50 C:\Users\Edu\AppData\Local\Temp\IXP001.TMP\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 130 196 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9672 0 0
2
45219.3 2
0
13 Logic Switch~
5 130 160 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 A2
-6 -27 8 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7876 0 0
2
45219.3 1
0
13 Logic Switch~
5 131 230 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6369 0 0
2
45219.3 0
0
5 4049~
219 183 137 0 2 22
0 3 2
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 2 0
1 U
9172 0 0
2
45219.3 0
0
5 4049~
219 384 325 0 2 22
0 12 8
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 2 0
1 U
7100 0 0
2
45219.3 3
0
5 4049~
219 385 358 0 2 22
0 11 7
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 2 0
1 U
3820 0 0
2
45219.3 2
0
5 4049~
219 387 393 0 2 22
0 10 6
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 1 0
1 U
7678 0 0
2
45219.3 1
0
5 4049~
219 384 290 0 2 22
0 13 9
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 1 0
1 U
961 0 0
2
45219.3 0
0
14 Logic Display~
6 567 128 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3178 0 0
2
45219.3 3
0
14 Logic Display~
6 619 128 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3409 0 0
2
45219.3 2
0
14 Logic Display~
6 594 128 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3951 0 0
2
45219.3 1
0
14 Logic Display~
6 645 127 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8885 0 0
2
45219.3 0
0
5 4049~
219 382 250 0 2 22
0 18 14
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 1 0
1 U
3780 0 0
2
45219.3 0
0
5 4049~
219 380 215 0 2 22
0 19 15
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 1 0
1 U
9265 0 0
2
45219.3 0
0
5 4049~
219 379 182 0 2 22
0 20 16
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 1 0
1 U
9442 0 0
2
45219.3 0
0
5 4049~
219 379 147 0 2 22
0 21 17
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
9424 0 0
2
45219.3 0
0
14 Logic Display~
6 490 129 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9968 0 0
2
45219.3 3
0
14 Logic Display~
6 515 129 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9281 0 0
2
45219.3 2
0
14 Logic Display~
6 541 128 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 1 0 0
1 L
8464 0 0
2
45219.3 1
0
14 Logic Display~
6 463 129 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7168 0 0
2
45219.3 0
0
7 74LS139
118 261 200 0 14 29
0 5 4 2 5 4 3 21 20 19
18 13 12 11 10
0
0 0 4848 0
7 74LS139
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 0
65 0 0 0 0 0 0 0
1 U
3171 0 0
2
45219.3 0
0
23
2 3 2 0 0 8336 0 4 21 0 0 4
204 137
224 137
224 200
223 200
0 1 3 0 0 4096 0 0 4 7 0 3
152 160
152 137
168 137
0 5 4 0 0 4096 0 0 21 5 0 3
215 207
215 227
229 227
0 4 5 0 0 8192 0 0 21 6 0 3
205 196
205 218
229 218
1 2 4 0 0 8320 0 3 21 0 0 5
143 230
143 207
215 207
215 191
229 191
1 1 5 0 0 4224 0 1 21 0 0 4
142 196
205 196
205 182
229 182
1 6 3 0 0 8320 0 2 21 0 0 4
142 160
152 160
152 236
223 236
1 2 6 0 0 4224 0 12 7 0 0 3
645 145
645 393
408 393
1 2 7 0 0 8320 0 10 6 0 0 3
619 146
619 358
406 358
1 2 8 0 0 8320 0 11 5 0 0 3
594 146
594 325
405 325
1 2 9 0 0 8320 0 9 8 0 0 3
567 146
567 290
405 290
14 1 10 0 0 8320 0 21 7 0 0 4
299 236
318 236
318 393
372 393
13 1 11 0 0 8320 0 21 6 0 0 4
299 227
326 227
326 358
370 358
12 1 12 0 0 8320 0 21 5 0 0 4
299 218
337 218
337 325
369 325
11 1 13 0 0 8320 0 21 8 0 0 4
299 209
346 209
346 290
369 290
2 1 14 0 0 4224 0 13 19 0 0 3
403 250
541 250
541 146
2 1 15 0 0 4224 0 14 18 0 0 3
401 215
515 215
515 147
2 1 16 0 0 4224 0 15 17 0 0 3
400 182
490 182
490 147
2 1 17 0 0 4224 0 16 20 0 0 2
400 147
463 147
10 1 18 0 0 4224 0 21 13 0 0 4
299 200
353 200
353 250
367 250
9 1 19 0 0 4224 0 21 14 0 0 4
299 191
362 191
362 215
365 215
8 1 20 0 0 4224 0 21 15 0 0 2
299 182
364 182
7 1 21 0 0 4224 0 21 16 0 0 4
299 173
361 173
361 147
364 147
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
