CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 30 120 10
225 411 1183 887
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
28 D:\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.500000 0.500000
225 411 1583 1134
42991634 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 107 561 0 1 11
0 33
0
0 0 21360 0
2 0V
-31 -1 -17 7
5 NUM15
-47 -13 -12 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
45373.4 0
0
13 Logic Switch~
5 105 538 0 1 11
0 29
0
0 0 21360 0
2 0V
-31 -1 -17 7
5 NUM14
-47 -13 -12 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
45373.4 1
0
13 Logic Switch~
5 106 516 0 1 11
0 28
0
0 0 21360 0
2 0V
-31 -1 -17 7
5 NUM13
-47 -13 -12 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
45373.4 2
0
13 Logic Switch~
5 107 493 0 1 11
0 27
0
0 0 21360 0
2 0V
-31 -1 -17 7
5 NUM12
-47 -13 -12 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
45373.4 3
0
13 Logic Switch~
5 107 471 0 1 11
0 26
0
0 0 21360 0
2 0V
-31 -1 -17 7
5 NUM11
-47 -13 -12 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
45373.4 4
0
13 Logic Switch~
5 99 238 0 1 11
0 34
0
0 0 21360 0
2 0V
-31 -1 -17 7
4 NUM1
-44 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
45373.4 5
0
13 Logic Switch~
5 99 259 0 1 11
0 32
0
0 0 21360 0
2 0V
-31 -1 -17 7
4 NUM2
-44 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
45373.4 6
0
13 Logic Switch~
5 101 284 0 1 11
0 31
0
0 0 21360 0
2 0V
-31 -1 -17 7
4 NUM3
-44 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
45373.4 7
0
13 Logic Switch~
5 102 309 0 1 11
0 30
0
0 0 21360 0
2 0V
-31 -1 -17 7
4 NUM4
-44 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
45373.4 8
0
13 Logic Switch~
5 102 334 0 1 11
0 22
0
0 0 21360 0
2 0V
-31 -1 -17 7
4 NUM5
-44 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
45373.4 9
0
13 Logic Switch~
5 102 356 0 1 11
0 21
0
0 0 21360 0
2 0V
-31 -1 -17 7
4 NUM6
-44 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
45373.4 10
0
13 Logic Switch~
5 103 380 0 1 11
0 20
0
0 0 21360 0
2 0V
-31 -1 -17 7
4 NUM7
-44 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
45373.4 11
0
13 Logic Switch~
5 104 404 0 1 11
0 23
0
0 0 21360 0
2 0V
-31 -1 -17 7
4 NUM8
-44 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
45373.4 12
0
13 Logic Switch~
5 106 427 0 1 11
0 24
0
0 0 21360 0
2 0V
-31 -1 -17 7
4 NUM9
-44 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4597 0 0
2
45373.4 13
0
13 Logic Switch~
5 107 450 0 1 11
0 25
0
0 0 21360 0
2 0V
-31 -1 -17 7
5 NUM10
-47 -13 -12 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3835 0 0
2
45373.4 14
0
12 DEC_BCH_7SEG
94 706 312 0 11 23
0 12 11 10 9 35 36 37 38 39
40 41
12 DEC_BCH_7SEG
1 0 4752 0
0
2 U2
-7 -55 7 -47
0
0
0
0
0
0
23

0 1 2 3 4 10 11 12 13 14
15 16 1 2 3 4 10 11 12 13
14 15 16 0
0 0 0 0 1 0 0 0
1 U
3670 0 0
2
45373.4 15
0
11 COD_HEX_BCH
94 306 384 0 19 39
0 34 32 31 30 22 21 20 23 24
25 26 27 28 29 33 9 10 11 12
11 COD_HEX_BCH
2 0 4784 0
0
2 U1
9 -86 23 -78
0
0
0
0
0
0
39

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 27 28 29 30
1 2 3 4 5 6 7 8 9 10
11 12 13 14 15 27 28 29 30 0
0 0 0 0 1 0 0 0
1 U
5616 0 0
2
45373.4 16
0
9 CC 7-Seg~
183 845 223 0 18 19
10 41 40 39 38 37 36 35 127 128
1 1 1 1 1 1 0 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9323 0 0
2
45373.4 17
0
26
16 4 9 0 0 4224 0 17 16 0 0 4
355 354
650 354
650 312
673 312
17 3 10 0 0 4224 0 17 16 0 0 4
355 345
655 345
655 303
673 303
18 2 11 0 0 4224 0 17 16 0 0 4
355 336
660 336
660 294
673 294
19 1 12 0 0 4224 0 17 16 0 0 4
355 327
665 327
665 285
673 285
1 7 20 0 0 12416 0 12 17 0 0 4
115 380
130 380
130 381
289 381
1 6 21 0 0 4224 0 11 17 0 0 4
114 356
243 356
243 372
289 372
1 5 22 0 0 4224 0 10 17 0 0 4
114 334
250 334
250 363
289 363
1 8 23 0 0 4224 0 13 17 0 0 4
116 404
237 404
237 390
289 390
1 9 24 0 0 4224 0 14 17 0 0 4
118 427
240 427
240 399
289 399
1 10 25 0 0 4224 0 15 17 0 0 4
119 450
245 450
245 408
289 408
1 11 26 0 0 4224 0 5 17 0 0 4
119 471
250 471
250 417
289 417
1 12 27 0 0 4224 0 4 17 0 0 4
119 493
255 493
255 426
289 426
1 13 28 0 0 4224 0 3 17 0 0 4
118 516
260 516
260 435
289 435
1 14 29 0 0 4224 0 2 17 0 0 4
117 538
265 538
265 444
289 444
1 4 30 0 0 4224 0 9 17 0 0 4
114 309
255 309
255 354
289 354
1 3 31 0 0 4224 0 8 17 0 0 4
113 284
260 284
260 345
289 345
1 2 32 0 0 4224 0 7 17 0 0 4
111 259
265 259
265 336
289 336
1 15 33 0 0 4224 0 1 17 0 0 4
119 561
270 561
270 453
289 453
1 1 34 0 0 4224 0 6 17 0 0 4
111 238
270 238
270 327
289 327
5 7 35 0 0 4224 0 16 18 0 0 3
739 339
860 339
860 259
6 6 36 0 0 4224 0 16 18 0 0 3
739 330
854 330
854 259
7 5 37 0 0 4224 0 16 18 0 0 3
739 321
848 321
848 259
8 4 38 0 0 4224 0 16 18 0 0 3
739 312
842 312
842 259
9 3 39 0 0 4224 0 16 18 0 0 3
739 303
836 303
836 259
10 2 40 0 0 4224 0 16 18 0 0 3
739 294
830 294
830 259
11 1 41 0 0 4224 0 16 18 0 0 3
739 285
824 285
824 259
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
