CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 30 30 110 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 1
20 Package,Description,
48 C:\Program Files (x86)\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 114 246 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
317 0 0
2
45226.3 0
0
13 Logic Switch~
5 114 212 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3108 0 0
2
45226.3 0
0
13 Logic Switch~
5 113 178 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4299 0 0
2
45226.3 0
0
13 Logic Switch~
5 113 143 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9672 0 0
2
45226.3 0
0
5 4049~
219 612 315 0 2 22
0 4 7
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 4 0
1 U
7876 0 0
2
45226.3 0
0
5 4049~
219 609 281 0 2 22
0 2 8
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 3 0
1 U
6369 0 0
2
45226.3 0
0
5 4049~
219 608 248 0 2 22
0 6 9
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
9172 0 0
2
45226.3 0
0
5 4049~
219 602 216 0 2 22
0 5 10
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
7100 0 0
2
45226.3 0
0
5 4049~
219 597 185 0 2 22
0 4 11
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
3820 0 0
2
45226.3 0
0
5 4049~
219 596 155 0 2 22
0 3 12
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
7678 0 0
2
45226.3 0
0
5 4049~
219 592 123 0 2 22
0 2 13
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
961 0 0
2
45226.3 0
0
14 Logic Display~
6 748 261 0 1 2
10 16
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3178 0 0
2
45226.3 5
0
14 Logic Display~
6 751 200 0 1 2
10 15
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3409 0 0
2
45226.3 4
0
14 Logic Display~
6 751 138 0 1 2
10 14
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L3
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3951 0 0
2
45226.3 3
0
8 3-In OR~
219 666 265 0 4 22
0 9 8 7 16
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 1 0
1 U
8885 0 0
2
45226.3 2
0
5 4071~
219 664 204 0 3 22
0 11 10 15
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
3780 0 0
2
45226.3 1
0
5 4071~
219 663 142 0 3 22
0 13 12 14
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
9265 0 0
2
45226.3 0
0
6 74LS42
101 306 188 0 14 29
0 20 19 18 17 21 22 23 6 5
24 2 3 4 25
0
0 0 4848 0
6 74LS42
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
106 %D [%16bi %8bi %1i %2i %3i %4i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 11 10 9 7 6
5 4 3 2 1 12 13 14 15 11
10 9 7 6 5 4 3 2 1 0
65 0 0 512 0 0 0 0
1 U
9442 0 0
2
45226.3 0
0
21
0 1 2 0 0 4096 0 0 11 6 0 3
529 281
529 123
577 123
12 1 3 0 0 4224 0 18 10 0 0 4
344 215
538 215
538 155
581 155
0 1 4 0 0 4112 0 0 9 7 0 3
568 315
568 185
582 185
9 1 5 0 0 4224 0 18 8 0 0 4
344 188
546 188
546 216
587 216
8 1 6 0 0 12416 0 18 7 0 0 4
344 179
436 179
436 248
593 248
11 1 2 0 0 12416 0 18 6 0 0 4
344 206
426 206
426 281
594 281
13 1 4 0 0 12416 0 18 5 0 0 4
344 224
419 224
419 315
597 315
2 3 7 0 0 4224 0 5 15 0 0 3
633 315
633 274
653 274
2 2 8 0 0 8320 0 6 15 0 0 3
630 281
630 265
654 265
2 1 9 0 0 8320 0 7 15 0 0 3
629 248
629 256
653 256
2 2 10 0 0 4224 0 8 16 0 0 4
623 216
652 216
652 213
651 213
2 1 11 0 0 8320 0 9 16 0 0 3
618 185
618 195
651 195
2 2 12 0 0 8320 0 10 17 0 0 3
617 155
617 151
650 151
2 1 13 0 0 8320 0 11 17 0 0 3
613 123
613 133
650 133
3 1 14 0 0 4224 0 17 14 0 0 2
696 142
735 142
3 1 15 0 0 4224 0 16 13 0 0 2
697 204
735 204
1 4 16 0 0 4224 0 12 15 0 0 2
732 265
699 265
1 4 17 0 0 4224 0 1 18 0 0 4
126 246
266 246
266 233
274 233
1 3 18 0 0 4224 0 2 18 0 0 4
126 212
250 212
250 224
274 224
1 2 19 0 0 4224 0 3 18 0 0 4
125 178
261 178
261 215
274 215
1 1 20 0 0 4224 0 4 18 0 0 4
125 143
266 143
266 206
274 206
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
