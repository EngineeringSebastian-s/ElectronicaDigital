CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
50 C:\Users\Edu\AppData\Local\Temp\IXP001.TMP\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
35
13 Logic Switch~
5 753 195 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 C2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9442 0 0
2
5.90094e-315 5.32571e-315
0
13 Logic Switch~
5 788 195 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 D2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9424 0 0
2
5.90094e-315 5.30499e-315
0
13 Logic Switch~
5 719 196 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 B2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9968 0 0
2
5.90094e-315 5.26354e-315
0
13 Logic Switch~
5 684 196 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 A2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9281 0 0
2
5.90094e-315 0
0
13 Logic Switch~
5 168 198 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
1 C
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8464 0 0
2
5.90094e-315 5.26354e-315
0
13 Logic Switch~
5 203 198 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
1 D
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7168 0 0
2
5.90094e-315 0
0
13 Logic Switch~
5 134 199 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3171 0 0
2
5.90094e-315 0
0
13 Logic Switch~
5 99 199 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4139 0 0
2
5.90094e-315 0
0
5 4081~
219 910 237 0 3 22
0 8 16 13
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 9 0
1 U
6435 0 0
2
5.90094e-315 5.41896e-315
0
14 Logic Display~
6 1222 286 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5283 0 0
2
5.90094e-315 5.41378e-315
0
5 4073~
219 989 312 0 4 22
0 10 7 9 4
0
0 0 608 0
4 4073
-7 -24 21 -16
4 U10C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 13 0
1 U
6874 0 0
2
5.90094e-315 5.4086e-315
0
8 4-In OR~
219 1109 381 0 5 22
0 13 4 12 5 11
0
0 0 608 0
4 4072
-14 -24 14 -16
3 U5B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 7 0
1 U
5305 0 0
2
5.90094e-315 5.40342e-315
0
5 4073~
219 993 397 0 4 22
0 2 15 9 12
0
0 0 608 0
4 4073
-7 -24 21 -16
4 U10B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 13 0
1 U
34 0 0
2
5.90094e-315 5.39824e-315
0
5 4073~
219 991 508 0 4 22
0 3 10 14 5
0
0 0 608 0
4 4073
-7 -24 21 -16
4 U10A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 13 0
1 U
969 0 0
2
5.90094e-315 5.39306e-315
0
5 4069~
219 838 244 0 2 22
0 9 16
0
0 0 608 0
4 4069
-7 -24 21 -16
3 U8D
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 4 12 0
1 U
8402 0 0
2
5.90094e-315 5.38788e-315
0
5 4069~
219 834 399 0 2 22
0 7 15
0
0 0 608 0
4 4069
-7 -24 21 -16
3 U8C
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 3 12 0
1 U
3751 0 0
2
5.90094e-315 5.37752e-315
0
5 4069~
219 834 466 0 2 22
0 8 3
0
0 0 608 0
4 4069
-7 -24 21 -16
3 U8B
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 2 12 0
1 U
4292 0 0
2
5.90094e-315 5.36716e-315
0
5 4069~
219 834 523 0 2 22
0 7 14
0
0 0 608 0
4 4069
-7 -24 21 -16
3 U8A
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 1 12 0
1 U
6118 0 0
2
5.90094e-315 5.3568e-315
0
5 4069~
219 834 355 0 2 22
0 8 2
0
0 0 608 0
4 4069
-7 -24 21 -16
3 U3F
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 6 10 0
1 U
34 0 0
2
5.90094e-315 5.34643e-315
0
5 4069~
219 249 526 0 2 22
0 18 32
0
0 0 608 0
4 4069
-7 -24 21 -16
3 U6E
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 5 8 0
1 U
6357 0 0
2
5.90094e-315 0
0
5 4069~
219 250 469 0 2 22
0 19 33
0
0 0 608 0
4 4069
-7 -24 21 -16
3 U6D
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 4 8 0
1 U
319 0 0
2
5.90094e-315 0
0
5 4069~
219 250 402 0 2 22
0 18 34
0
0 0 608 0
4 4069
-7 -24 21 -16
3 U6C
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 3 8 0
1 U
3976 0 0
2
5.90094e-315 0
0
5 4069~
219 250 365 0 2 22
0 19 35
0
0 0 608 0
4 4069
-7 -24 21 -16
3 U6B
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 2 8 0
1 U
7634 0 0
2
5.90094e-315 0
0
5 4069~
219 250 247 0 2 22
0 20 36
0
0 0 608 0
4 4069
-7 -24 21 -16
3 U6A
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 1 8 0
1 U
523 0 0
2
5.90094e-315 0
0
5 4071~
219 582 378 0 3 22
0 23 24 22
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 6 0
1 U
6748 0 0
2
5.90094e-315 0
0
5 4071~
219 504 459 0 3 22
0 26 25 24
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
6901 0 0
2
5.90094e-315 0
0
5 4071~
219 503 292 0 3 22
0 28 27 23
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
842 0 0
2
5.90094e-315 0
0
5 4081~
219 402 511 0 3 22
0 31 32 25
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
3277 0 0
2
5.90094e-315 0
0
5 4081~
219 332 486 0 3 22
0 33 21 31
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
4212 0 0
2
5.90094e-315 0
0
5 4081~
219 402 417 0 3 22
0 30 20 26
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
4720 0 0
2
5.90094e-315 0
0
5 4081~
219 401 331 0 3 22
0 29 20 27
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
5551 0 0
2
5.90094e-315 0
0
5 4081~
219 330 391 0 3 22
0 35 34 30
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
6986 0 0
2
5.90094e-315 0
0
5 4081~
219 329 312 0 3 22
0 21 18 29
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
8745 0 0
2
5.90094e-315 0
0
5 4081~
219 325 240 0 3 22
0 19 36 28
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
9592 0 0
2
5.90094e-315 0
0
14 Logic Display~
6 637 289 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8748 0 0
2
5.90094e-315 0
0
49
2 1 2 0 0 12416 0 19 13 0 0 5
855 355
883 355
883 381
969 381
969 388
2 1 3 0 0 4224 0 17 14 0 0 4
855 466
959 466
959 499
967 499
4 2 4 0 0 8320 0 11 12 0 0 4
1010 312
1067 312
1067 377
1092 377
4 4 5 0 0 8320 0 12 14 0 0 4
1092 395
1083 395
1083 508
1012 508
0 0 6 0 0 0 0 0 0 0 0 2
788 444
788 444
0 1 7 0 0 4096 0 0 16 20 0 2
753 399
819 399
0 1 8 0 0 4096 0 0 19 22 0 2
684 355
819 355
0 3 9 0 0 4096 0 0 11 19 0 3
788 328
965 328
965 321
0 2 7 0 0 4096 0 0 11 20 0 3
753 310
965 310
965 312
0 1 10 0 0 4096 0 0 11 21 0 3
719 282
965 282
965 303
0 1 9 0 0 0 0 0 15 19 0 2
788 244
823 244
0 1 8 0 0 4096 0 0 9 22 0 2
684 228
886 228
5 1 11 0 0 4224 0 12 10 0 0 3
1142 381
1222 381
1222 304
4 3 12 0 0 4224 0 13 12 0 0 4
1014 397
1067 397
1067 386
1092 386
3 1 13 0 0 4224 0 9 12 0 0 4
931 237
1085 237
1085 368
1092 368
2 3 14 0 0 4224 0 18 14 0 0 4
855 523
956 523
956 517
967 517
2 2 15 0 0 12416 0 16 13 0 0 4
855 399
883 399
883 397
969 397
2 2 16 0 0 4224 0 15 9 0 0 4
859 244
877 244
877 246
886 246
1 3 9 0 0 4224 0 2 13 0 0 4
788 207
788 435
969 435
969 406
1 1 7 0 0 4224 0 1 18 0 0 3
753 207
753 523
819 523
1 2 10 0 0 4224 0 3 14 0 0 5
719 208
719 491
893 491
893 508
967 508
1 1 8 0 0 4224 0 4 17 0 0 3
684 208
684 466
819 466
0 0 17 0 0 0 0 0 0 0 0 2
203 447
203 447
0 1 18 0 0 4096 0 0 22 47 0 2
168 402
235 402
0 1 19 0 0 4096 0 0 23 49 0 2
99 365
235 365
0 2 20 0 0 4096 0 0 31 46 0 2
203 340
377 340
0 2 18 0 0 4096 0 0 33 47 0 2
168 321
305 321
0 1 21 0 0 4096 0 0 33 48 0 2
134 303
305 303
0 1 20 0 0 0 0 0 24 46 0 2
203 247
235 247
0 1 19 0 0 4096 0 0 34 49 0 2
99 231
301 231
3 1 22 0 0 12416 0 25 35 0 0 4
615 378
615 377
637 377
637 307
3 1 23 0 0 8320 0 27 25 0 0 5
536 292
560 292
560 368
569 368
569 369
3 2 24 0 0 12416 0 26 25 0 0 6
537 459
537 460
560 460
560 386
569 386
569 387
3 2 25 0 0 4224 0 28 26 0 0 5
423 511
482 511
482 469
491 469
491 468
3 1 26 0 0 4224 0 30 26 0 0 5
423 417
482 417
482 451
491 451
491 450
3 2 27 0 0 4224 0 31 27 0 0 4
422 331
482 331
482 301
490 301
3 1 28 0 0 4224 0 34 27 0 0 4
346 240
482 240
482 283
490 283
3 1 29 0 0 4224 0 33 31 0 0 4
350 312
367 312
367 322
377 322
3 1 30 0 0 4224 0 32 30 0 0 4
351 391
369 391
369 408
378 408
3 1 31 0 0 8320 0 29 28 0 0 5
353 486
353 485
371 485
371 502
378 502
2 2 32 0 0 4224 0 20 28 0 0 4
270 526
371 526
371 520
378 520
2 1 33 0 0 4224 0 21 29 0 0 5
271 469
301 469
301 476
308 476
308 477
2 2 34 0 0 4224 0 22 32 0 0 4
271 402
298 402
298 400
306 400
2 1 35 0 0 4224 0 23 32 0 0 4
271 365
298 365
298 382
306 382
2 2 36 0 0 4224 0 24 34 0 0 4
271 247
292 247
292 249
301 249
1 2 20 0 0 4224 0 6 30 0 0 3
203 210
203 426
378 426
1 1 18 0 0 4224 0 5 20 0 0 3
168 210
168 526
234 526
1 2 21 0 0 4224 0 7 29 0 0 4
134 211
134 494
308 494
308 495
1 1 19 0 0 4224 0 8 21 0 0 3
99 211
99 469
235 469
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
129 103 246 127
139 111 235 127
12 Dos entradas
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
702 105 827 129
712 113 816 129
13 Tres entradas
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
234 104 391 128
244 112 380 128
17 A~D + BCD + ~A~CD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
381 104 458 128
391 112 447 128
7 + ~AB~C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
964 104 1041 128
974 112 1030 128
7 + ~AB~C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
815 104 972 128
825 112 961 128
17 A~D + BCD + ~A~CD
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
