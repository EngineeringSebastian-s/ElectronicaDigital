CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 130 30 150 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
50 C:\Users\Edu\AppData\Local\Temp\IXP000.TMP\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1702 537
9961490 0
0
6 Title:
5 Name:
0
0
0
30
7 Ground~
168 5 314 0 1 3
0 15
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 0 0 0 0
3 GND
3409 0 0
2
45177.3 0
0
11 Multimeter~
205 125 688 0 21 21
0 2 16 17 3 0 0 0 0 0
32 54 46 53 56 50 32 32 0 0
4 73
0
0 0 16464 90
6 1.000u
-21 -19 21 -11
3 MM0
-11 -29 10 -21
0
0
31 R1%D %1 %2 1E-9
%D %4 %2 DC %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
73 0 0 0 0 0 0 0
1 I
3951 0 0
2
45177.3 0
0
9 Resistor~
219 449 753 0 2 5
0 6 3
0
0 0 880 90
1 4
14 0 21 8
3 R28
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
8885 0 0
2
45177.3 0
0
9 Resistor~
219 359 806 0 2 5
0 2 6
0
0 0 880 0
1 8
-4 -14 3 -6
3 R27
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3780 0 0
2
45177.3 0
0
9 Resistor~
219 362 697 0 2 5
0 5 4
0
0 0 880 0
2 12
-7 -14 7 -6
3 R26
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9265 0 0
2
45177.3 0
0
9 Resistor~
219 510 697 0 2 5
0 4 6
0
0 0 880 0
2 12
-7 -14 7 -6
3 R25
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9442 0 0
2
45177.3 0
0
9 Resistor~
219 508 617 0 2 5
0 3 6
0
0 0 880 0
1 6
-4 -14 3 -6
3 R24
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9424 0 0
2
45177.3 0
0
9 Resistor~
219 263 756 0 2 5
0 2 5
0
0 0 880 90
1 2
14 0 21 8
3 R23
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9968 0 0
2
45177.3 0
0
9 Resistor~
219 264 653 0 2 5
0 5 3
0
0 0 880 90
2 24
11 0 25 8
3 R22
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9281 0 0
2
45177.3 0
0
9 Resistor~
219 530 458 0 2 5
0 10 7
0
0 0 880 0
2 1k
-7 -14 7 -6
3 R21
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
8464 0 0
2
45177.3 0
0
9 Resistor~
219 370 458 0 2 5
0 9 10
0
0 0 880 0
2 1k
-7 -14 7 -6
3 R20
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7168 0 0
2
45177.3 0
0
9 Resistor~
219 337 361 0 2 5
0 11 12
0
0 0 880 90
2 1k
11 0 25 8
3 R19
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3171 0 0
2
45177.3 0
0
9 Resistor~
219 314 323 0 2 5
0 9 12
0
0 0 880 0
2 1k
-7 -14 7 -6
3 R18
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
4139 0 0
2
45177.3 0
0
9 Resistor~
219 311 260 0 2 5
0 9 12
0
0 0 880 0
2 1k
-7 -14 7 -6
3 R17
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
6435 0 0
2
45177.3 0
0
9 Resistor~
219 649 246 0 2 5
0 13 8
0
0 0 880 90
2 1k
11 0 25 8
3 R16
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
5283 0 0
2
45177.3 0
0
9 Resistor~
219 678 331 0 2 5
0 8 7
0
0 0 880 0
2 1k
-7 -14 7 -6
3 R15
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
6874 0 0
2
45177.3 0
0
9 Resistor~
219 286 394 0 2 5
0 9 11
0
0 0 880 0
2 1k
-7 -14 7 -6
3 R14
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
5305 0 0
2
45177.3 0
0
9 Resistor~
219 211 296 0 2 5
0 9 14
0
0 0 880 90
2 1k
11 0 25 8
3 R13
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
34 0 0
2
45177.3 0
0
9 Resistor~
219 878 306 0 2 5
0 7 13
0
0 0 880 90
2 1k
11 0 25 8
3 R12
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
969 0 0
2
45177.3 0
0
9 Resistor~
219 390 310 0 2 5
0 11 12
0
0 0 880 90
2 1k
11 0 25 8
3 R11
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
8402 0 0
2
45177.3 0
0
9 Resistor~
219 957 293 0 2 5
0 7 13
0
0 0 880 90
2 1k
11 0 25 8
3 R10
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3751 0 0
2
45177.3 0
0
9 Resistor~
219 802 296 0 2 5
0 7 13
0
0 0 880 90
2 1k
8 0 22 8
2 R9
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
4292 0 0
2
45177.3 0
0
9 Resistor~
219 801 401 0 2 5
0 7 7
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
6118 0 0
2
45177.3 0
0
9 Resistor~
219 714 217 0 2 5
0 8 13
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
34 0 0
2
45177.3 0
0
9 Resistor~
219 586 293 0 2 5
0 8 13
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
6357 0 0
2
45177.3 0
0
9 Resistor~
219 586 390 0 2 5
0 8 7
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
319 0 0
2
45177.3 0
0
9 Resistor~
219 436 390 0 2 5
0 11 8
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3976 0 0
2
45177.3 0
0
9 Resistor~
219 489 296 0 2 5
0 8 8
0
0 0 880 90
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7634 0 0
2
45177.3 0
0
9 Resistor~
219 432 217 0 2 5
0 12 8
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
523 0 0
2
45177.3 0
0
9 Resistor~
219 318 219 0 2 5
0 14 12
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
6748 0 0
2
45177.3 0
0
49
1 0 2 0 0 8320 0 2 0 0 4 4
142 719
183 719
183 806
263 806
4 0 3 0 0 12288 0 2 0 0 12 4
142 669
185 669
185 617
264 617
0 1 4 0 0 4096 0 0 6 7 0 2
449 697
492 697
1 1 2 0 0 16 0 8 4 0 0 3
263 774
263 806
341 806
0 2 5 0 0 4096 0 0 8 6 0 3
264 697
264 738
263 738
1 1 5 0 0 8320 0 9 5 0 0 3
264 671
264 697
344 697
2 0 4 0 0 4224 0 5 0 0 0 3
380 697
449 697
449 690
1 0 6 0 0 4096 0 3 0 0 11 2
449 771
449 806
2 0 6 0 0 0 0 6 0 0 11 2
528 697
558 697
0 2 3 0 0 4096 0 0 3 12 0 2
449 617
449 735
2 2 6 0 0 8320 0 7 4 0 0 4
526 617
558 617
558 806
377 806
2 1 3 0 0 8320 0 9 7 0 0 3
264 635
264 617
490 617
0 0 7 0 0 4096 0 0 0 16 46 4
774 458
952 458
952 401
957 401
0 0 8 0 0 8192 0 0 0 43 48 3
560 296
546 296
546 217
0 0 9 0 0 4096 0 0 0 29 26 3
211 346
286 346
286 323
2 0 7 0 0 4224 0 10 0 0 42 4
548 458
774 458
774 401
779 401
2 1 10 0 0 4224 0 11 10 0 0 2
388 458
512 458
0 1 9 0 0 8320 0 0 11 29 0 3
211 394
211 458
352 458
1 0 11 0 0 4096 0 12 0 0 28 2
337 379
337 394
0 2 12 0 0 8192 0 0 12 27 0 3
340 319
337 319
337 343
0 0 13 0 0 4096 0 0 0 47 23 2
957 238
752 238
0 0 7 0 0 0 0 0 0 46 35 2
957 344
878 344
0 0 13 0 0 0 0 0 0 47 44 2
752 217
752 274
0 0 7 0 0 0 0 0 0 31 42 2
715 331
715 390
0 0 12 0 0 4096 0 0 0 27 38 2
340 274
390 274
1 1 9 0 0 0 0 13 14 0 0 4
296 323
285 323
285 260
293 260
2 2 12 0 0 8192 0 14 13 0 0 4
329 260
340 260
340 323
332 323
2 0 11 0 0 4224 0 17 0 0 37 4
304 394
385 394
385 390
390 390
1 1 9 0 0 0 0 18 17 0 0 3
211 314
211 394
268 394
2 1 14 0 0 8320 0 18 30 0 0 3
211 278
211 219
300 219
2 0 7 0 0 0 0 16 0 0 45 4
696 331
774 331
774 332
779 332
0 1 8 0 0 4096 0 0 16 43 0 2
560 331
660 331
2 0 8 0 0 0 0 15 0 0 48 4
649 228
649 222
650 222
650 217
1 0 13 0 0 0 0 15 0 0 44 3
649 264
649 274
650 274
1 0 7 0 0 0 0 19 0 0 46 2
878 324
878 401
0 2 13 0 0 0 0 0 19 44 0 3
802 274
878 274
878 288
1 1 11 0 0 0 0 20 27 0 0 3
390 328
390 390
418 390
2 0 12 0 0 4224 0 20 0 0 49 2
390 292
390 219
2 0 8 0 0 4096 0 27 0 0 43 2
454 390
560 390
2 0 8 0 0 0 0 28 0 0 48 2
489 278
489 217
0 1 8 0 0 0 0 0 28 43 0 3
560 329
489 329
489 314
2 0 7 0 0 0 0 26 0 0 45 3
604 390
779 390
779 401
1 1 8 0 0 0 0 25 26 0 0 4
568 293
560 293
560 390
568 390
2 2 13 0 0 0 0 22 25 0 0 5
802 278
802 274
612 274
612 293
604 293
1 1 7 0 0 0 0 23 22 0 0 5
783 401
779 401
779 322
802 322
802 314
1 2 7 0 0 0 0 21 23 0 0 3
957 311
957 401
819 401
2 2 13 0 0 4224 0 24 21 0 0 3
732 217
957 217
957 275
2 1 8 0 0 4224 0 29 24 0 0 2
450 217
696 217
2 1 12 0 0 0 0 30 29 0 0 4
336 219
406 219
406 217
414 217
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
