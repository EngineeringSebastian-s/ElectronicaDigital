CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 1
20 Package,Description,
48 C:\Program Files (x86)\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
50
13 Logic Switch~
5 99 340 0 1 11
0 47
0
0 0 21360 0
2 0V
-38 -1 -24 7
4 NUM1
-43 -13 -15 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3372 0 0
2
45226.5 0
0
13 Logic Switch~
5 97 211 0 1 11
0 51
0
0 0 21360 0
2 0V
-38 -1 -24 7
4 NUM5
-44 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3741 0 0
2
45226.5 1
0
13 Logic Switch~
5 97 241 0 1 11
0 50
0
0 0 21360 0
2 0V
-38 -1 -24 7
4 NUM4
-44 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5813 0 0
2
45226.5 2
0
13 Logic Switch~
5 98 275 0 1 11
0 49
0
0 0 21360 0
2 0V
-38 -1 -24 7
4 NUM3
-44 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3213 0 0
2
45226.5 3
0
13 Logic Switch~
5 98 305 0 1 11
0 48
0
0 0 21360 0
2 0V
-38 -1 -24 7
4 NUM2
-44 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3694 0 0
2
45226.5 4
0
13 Logic Switch~
5 96 146 0 1 11
0 53
0
0 0 21360 0
2 0V
-38 -1 -24 7
4 NUM7
-44 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4327 0 0
2
45226.5 5
0
13 Logic Switch~
5 96 176 0 1 11
0 52
0
0 0 21360 0
2 0V
-38 -1 -24 7
4 NUM6
-44 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8800 0 0
2
45226.5 6
0
13 Logic Switch~
5 95 112 0 1 11
0 54
0
0 0 21360 0
2 0V
-38 -1 -24 7
4 NUM8
-44 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3406 0 0
2
45226.5 7
0
13 Logic Switch~
5 95 82 0 1 11
0 55
0
0 0 21360 0
2 0V
-38 -1 -24 7
4 NUM9
-44 -13 -16 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6455 0 0
2
45226.5 8
0
6 74LS48
188 455 527 0 14 29
0 22 20 19 21 60 61 12 13 14
15 16 17 18 62
0
0 0 4848 0
7 74LS248
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9319 0 0
2
45226.5 24
0
5 4049~
219 381 528 0 2 22
0 24 19
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 4 0
1 U
3172 0 0
2
45226.5 23
0
5 4049~
219 381 483 0 2 22
0 25 20
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 4 0
1 U
38 0 0
2
45226.5 22
0
5 4049~
219 346 561 0 2 22
0 23 21
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 4 0
1 U
376 0 0
2
45226.5 21
0
5 4049~
219 347 461 0 2 22
0 26 22
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 4 0
1 U
6666 0 0
2
45226.5 20
0
5 74147
219 267 526 0 13 27
0 11 10 9 8 7 6 5 4 3
23 24 25 26
0
0 0 4848 0
5 74147
-18 -60 17 -52
2 U8
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
121 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
27

0 10 5 4 3 2 1 13 12 11
9 7 6 14 10 5 4 3 2 1
13 12 11 9 7 6 14 0
65 0 0 0 1 0 0 0
1 U
9365 0 0
2
45226.5 19
0
9 CC 7-Seg~
183 732 444 0 18 19
10 18 17 16 15 14 13 12 63 64
1 1 1 1 1 1 0 2 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3251 0 0
2
45226.5 18
0
14 NO PushButton~
191 110 490 0 2 5
0 10 2
0
0 0 4720 0
0
4 NUM8
-37 -10 -9 -2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
5481 0 0
2
45226.5 17
0
14 NO PushButton~
191 111 457 0 2 5
0 11 2
0
0 0 4720 0
0
4 NUM9
-37 -10 -9 -2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
7788 0 0
2
45226.5 16
0
14 NO PushButton~
191 109 516 0 2 5
0 9 2
0
0 0 4720 0
0
4 NUM7
-37 -10 -9 -2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
3273 0 0
2
45226.5 15
0
14 NO PushButton~
191 110 546 0 2 5
0 8 2
0
0 0 4720 0
0
4 NUM6
-37 -10 -9 -2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
3761 0 0
2
45226.5 14
0
14 NO PushButton~
191 108 636 0 2 5
0 5 2
0
0 0 4720 0
0
4 NUM3
-37 -10 -9 -2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
3226 0 0
2
45226.5 13
0
14 NO PushButton~
191 109 610 0 2 5
0 6 2
0
0 0 4720 0
0
4 NUM4
-37 -10 -9 -2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
4244 0 0
2
45226.5 12
0
14 NO PushButton~
191 108 580 0 2 5
0 7 2
0
0 0 4720 0
0
4 NUM5
-37 -10 -9 -2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
5225 0 0
2
45226.5 11
0
14 NO PushButton~
191 109 666 0 2 5
0 4 2
0
0 0 4720 0
0
4 NUM2
-37 -10 -9 -2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
768 0 0
2
45226.5 10
0
14 NO PushButton~
191 110 695 0 2 5
0 3 2
0
0 0 4720 0
0
4 NUM1
-36 -10 -8 -2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 0 0 0 0
1 S
5735 0 0
2
45226.5 9
0
7 Ground~
168 88 464 0 1 3
0 2
0
0 0 53360 270
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5881 0 0
2
45226.5 8
0
7 Ground~
168 87 497 0 1 3
0 2
0
0 0 53360 270
0
4 GND2
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3275 0 0
2
45226.5 7
0
7 Ground~
168 86 523 0 1 3
0 2
0
0 0 53360 270
0
4 GND3
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4203 0 0
2
45226.5 6
0
7 Ground~
168 87 553 0 1 3
0 2
0
0 0 53360 270
0
4 GND4
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3440 0 0
2
45226.5 5
0
7 Ground~
168 85 587 0 1 3
0 2
0
0 0 53360 270
0
4 GND5
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9102 0 0
2
45226.5 4
0
7 Ground~
168 86 617 0 1 3
0 2
0
0 0 53360 270
0
4 GND6
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5586 0 0
2
45226.5 3
0
7 Ground~
168 84 643 0 1 3
0 2
0
0 0 53360 270
0
4 GND7
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
525 0 0
2
45226.5 2
0
7 Ground~
168 86 673 0 1 3
0 2
0
0 0 53360 270
0
4 GND8
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6206 0 0
2
45226.5 1
0
7 Ground~
168 86 702 0 1 3
0 2
0
0 0 53360 270
0
4 GND9
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3418 0 0
2
45226.5 0
0
6 74LS48
188 484 150 0 14 29
0 37 35 34 36 65 66 27 28 29
30 31 32 33 67
0
0 0 4848 0
7 74LS248
-24 -60 25 -52
2 U7
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9312 0 0
2
5.90098e-315 0
0
5 4049~
219 410 151 0 2 22
0 57 34
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 4 0
1 U
7419 0 0
2
45226.5 9
0
5 4049~
219 410 106 0 2 22
0 58 35
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 4 0
1 U
472 0 0
2
45226.5 10
0
5 4049~
219 375 184 0 2 22
0 56 36
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 3 0
1 U
4714 0 0
2
45226.5 11
0
5 4049~
219 376 84 0 2 22
0 59 37
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
9386 0 0
2
45226.5 12
0
5 4049~
219 147 369 0 2 22
0 47 38
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 2 0
1 U
7610 0 0
2
45226.5 13
0
5 4049~
219 167 335 0 2 22
0 48 39
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 2 0
1 U
3482 0 0
2
45226.5 14
0
5 4049~
219 189 304 0 2 22
0 49 40
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 2 0
1 U
3608 0 0
2
45226.5 15
0
5 4049~
219 189 269 0 2 22
0 50 41
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 1 0
1 U
6397 0 0
2
45226.5 16
0
5 4049~
219 160 209 0 2 22
0 51 42
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 1 0
1 U
3967 0 0
2
45226.5 17
0
5 4049~
219 214 119 0 2 22
0 52 43
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 1 0
1 U
8621 0 0
2
45226.5 18
0
5 4049~
219 190 96 0 2 22
0 53 44
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 1 0
1 U
8901 0 0
2
45226.5 19
0
5 4049~
219 168 76 0 2 22
0 54 45
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 1 0
1 U
7385 0 0
2
45226.5 20
0
5 4049~
219 146 52 0 2 22
0 55 46
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
6519 0 0
2
45226.5 21
0
5 74147
219 300 142 0 13 27
0 46 45 44 43 42 41 40 39 38
56 57 58 59
0
0 0 4848 0
5 74147
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
121 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
27

0 10 5 4 3 2 1 13 12 11
9 7 6 14 10 5 4 3 2 1
13 12 11 9 7 6 14 0
65 0 0 0 1 0 0 0
1 U
552 0 0
2
45226.5 22
0
9 CC 7-Seg~
183 761 67 0 18 19
10 33 32 31 30 29 28 27 68 69
1 1 1 1 1 1 0 2 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5551 0 0
2
45226.5 23
0
66
1 2 2 0 0 16 0 34 25 0 0 2
93 703
93 703
1 2 2 0 0 4240 0 33 24 0 0 2
93 674
92 674
1 2 2 0 0 16 0 32 21 0 0 2
91 644
91 644
1 2 2 0 0 16 0 31 22 0 0 2
93 618
92 618
1 2 2 0 0 16 0 30 23 0 0 2
92 588
91 588
1 2 2 0 0 16 0 29 20 0 0 2
94 554
93 554
1 2 2 0 0 16 0 28 19 0 0 2
93 524
92 524
1 2 2 0 0 16 0 27 17 0 0 2
94 498
93 498
1 2 2 0 0 16 0 26 18 0 0 2
95 465
94 465
1 9 3 0 0 8336 0 25 15 0 0 4
127 703
228 703
228 562
229 562
1 8 4 0 0 8336 0 24 15 0 0 4
126 674
224 674
224 553
229 553
1 7 5 0 0 8336 0 21 15 0 0 4
125 644
219 644
219 544
229 544
1 6 6 0 0 4240 0 22 15 0 0 4
126 618
215 618
215 535
229 535
1 5 7 0 0 4240 0 23 15 0 0 4
125 588
209 588
209 526
229 526
1 4 8 0 0 4240 0 20 15 0 0 4
127 554
204 554
204 517
229 517
1 3 9 0 0 4240 0 19 15 0 0 4
126 524
200 524
200 508
229 508
1 2 10 0 0 4240 0 17 15 0 0 4
127 498
221 498
221 499
229 499
1 1 11 0 0 4240 0 18 15 0 0 4
128 465
221 465
221 490
229 490
7 7 12 0 0 4240 0 10 16 0 0 3
487 491
747 491
747 480
8 6 13 0 0 4240 0 10 16 0 0 3
487 500
741 500
741 480
9 5 14 0 0 4240 0 10 16 0 0 3
487 509
735 509
735 480
10 4 15 0 0 4240 0 10 16 0 0 3
487 518
729 518
729 480
11 3 16 0 0 4240 0 10 16 0 0 3
487 527
723 527
723 480
12 2 17 0 0 4240 0 10 16 0 0 3
487 536
717 536
717 480
13 1 18 0 0 4240 0 10 16 0 0 3
487 545
711 545
711 480
2 3 19 0 0 8336 0 11 10 0 0 4
402 528
406 528
406 509
423 509
2 2 20 0 0 12432 0 12 10 0 0 4
402 483
405 483
405 500
423 500
2 4 21 0 0 4240 0 13 10 0 0 4
367 561
413 561
413 518
423 518
2 1 22 0 0 8336 0 14 10 0 0 5
368 461
368 462
414 462
414 491
423 491
10 1 23 0 0 8336 0 15 13 0 0 4
305 535
320 535
320 561
331 561
11 1 24 0 0 12432 0 15 11 0 0 4
305 526
328 526
328 528
366 528
12 1 25 0 0 12432 0 15 12 0 0 4
305 517
328 517
328 483
366 483
13 1 26 0 0 8336 0 15 14 0 0 4
305 508
318 508
318 461
332 461
7 7 27 0 0 4224 0 35 50 0 0 3
516 114
776 114
776 103
8 6 28 0 0 4224 0 35 50 0 0 3
516 123
770 123
770 103
9 5 29 0 0 4224 0 35 50 0 0 3
516 132
764 132
764 103
10 4 30 0 0 4224 0 35 50 0 0 3
516 141
758 141
758 103
11 3 31 0 0 4224 0 35 50 0 0 3
516 150
752 150
752 103
12 2 32 0 0 4224 0 35 50 0 0 3
516 159
746 159
746 103
13 1 33 0 0 4224 0 35 50 0 0 3
516 168
740 168
740 103
2 3 34 0 0 8320 0 36 35 0 0 4
431 151
435 151
435 132
452 132
2 2 35 0 0 12416 0 37 35 0 0 4
431 106
434 106
434 123
452 123
2 4 36 0 0 4224 0 38 35 0 0 4
396 184
442 184
442 141
452 141
2 1 37 0 0 8320 0 39 35 0 0 5
397 84
397 85
443 85
443 114
452 114
2 9 38 0 0 8320 0 40 49 0 0 4
168 369
249 369
249 178
262 178
2 8 39 0 0 8320 0 41 49 0 0 4
188 335
244 335
244 169
262 169
2 7 40 0 0 8320 0 42 49 0 0 4
210 304
239 304
239 160
262 160
2 6 41 0 0 8320 0 43 49 0 0 4
210 269
223 269
223 151
262 151
2 5 42 0 0 8320 0 44 49 0 0 4
181 209
203 209
203 142
262 142
2 4 43 0 0 12416 0 45 49 0 0 4
235 119
241 119
241 133
262 133
2 3 44 0 0 4224 0 46 49 0 0 4
211 96
245 96
245 124
262 124
2 2 45 0 0 4224 0 47 49 0 0 4
189 76
253 76
253 115
262 115
2 1 46 0 0 4224 0 48 49 0 0 4
167 52
259 52
259 106
262 106
1 1 47 0 0 8320 0 1 40 0 0 4
111 340
121 340
121 369
132 369
1 1 48 0 0 8320 0 5 41 0 0 4
110 305
134 305
134 335
152 335
1 1 49 0 0 12416 0 4 42 0 0 4
110 275
141 275
141 304
174 304
1 1 50 0 0 4224 0 3 43 0 0 4
109 241
146 241
146 269
174 269
1 1 51 0 0 12416 0 2 44 0 0 4
109 211
120 211
120 209
145 209
1 1 52 0 0 8320 0 7 45 0 0 4
108 176
144 176
144 119
199 119
1 1 53 0 0 8320 0 6 46 0 0 4
108 146
135 146
135 96
175 96
1 1 54 0 0 8320 0 8 47 0 0 4
107 112
128 112
128 76
153 76
1 1 55 0 0 8320 0 9 48 0 0 4
107 82
119 82
119 52
131 52
10 1 56 0 0 8320 0 49 38 0 0 4
338 151
349 151
349 184
360 184
11 1 57 0 0 12416 0 49 36 0 0 4
338 142
357 142
357 151
395 151
12 1 58 0 0 12416 0 49 37 0 0 4
338 133
357 133
357 106
395 106
13 1 59 0 0 8320 0 49 39 0 0 4
338 124
347 124
347 84
361 84
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
