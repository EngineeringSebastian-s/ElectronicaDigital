CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 330 30 100 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
50 C:\Users\Edu\AppData\Local\Temp\IXP000.TMP\BOM.DAT
0 7
2 4 0.499308 0.500000
344 176 1702 537
9961490 0
0
6 Title:
5 Name:
0
0
0
18
11 Multimeter~
205 262 676 0 21 21
0 3 17 18 2 0 0 0 0 0
32 55 46 54 56 48 32 32 0 0
4 73
0
0 0 16464 90
6 1.000u
-21 -19 21 -11
3 MM5
-11 -29 10 -21
0
0
31 R1%D %1 %2 1E-9
%D %4 %2 DC %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
73 0 0 0 0 0 0 0
1 I
317 0 0
2
45174.3 0
0
11 Multimeter~
205 262 555 0 21 21
0 5 19 20 6 0 0 0 0 0
32 55 46 54 56 48 32 32 0 0
4 73
0
0 0 16464 90
6 1.000u
-21 -19 21 -11
3 MM4
-11 -29 10 -21
0
0
31 R1%D %1 %2 1E-9
%D %4 %2 DC %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
73 0 0 0 0 0 0 0
1 I
3108 0 0
2
45174.3 0
0
11 Multimeter~
205 262 432 0 21 21
0 9 21 22 10 0 0 0 0 0
32 55 46 54 56 52 32 32 0 0
4 73
0
0 0 16464 90
6 1.000u
-21 -19 21 -11
3 MM3
-11 -29 10 -21
0
0
31 R1%D %1 %2 1E-9
%D %4 %2 DC %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
73 0 0 0 0 0 0 0
1 I
4299 0 0
2
45174.3 0
0
7 Ground~
168 192 404 0 1 3
0 23
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 0 0 0 0
3 GND
9672 0 0
2
45174.3 0
0
11 Multimeter~
205 262 300 0 21 21
0 12 24 25 13 0 0 0 0 0
32 55 46 54 56 52 32 32 0 0
4 73
0
0 0 16464 90
6 1.000u
-21 -19 21 -11
3 MM0
-11 -29 10 -21
0
0
31 R1%D %1 %2 1E-9
%D %4 %2 DC %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
73 0 0 0 0 0 0 0
1 I
7876 0 0
2
45174.3 0
0
9 Resistor~
219 421 686 0 2 5
0 3 2
0
0 0 880 90
4 7.68
1 0 29 8
3 R13
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
6369 0 0
2
45174.3 1
0
9 Resistor~
219 421 565 0 2 5
0 7 4
0
0 0 880 90
4 3.68
1 0 29 8
3 R12
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9172 0 0
2
45174.3 3
0
9 Resistor~
219 384 611 0 2 5
0 5 7
0
0 0 880 0
1 1
-4 -14 3 -6
3 R11
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7100 0 0
2
45174.3 2
0
9 Resistor~
219 382 518 0 2 5
0 6 4
0
0 0 880 0
1 3
-4 -14 3 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3820 0 0
2
45174.3 1
0
9 Resistor~
219 382 395 0 2 5
0 10 8
0
0 0 880 0
1 3
-4 -14 3 -6
3 R10
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7678 0 0
2
45174.3 5
0
9 Resistor~
219 384 488 0 2 5
0 9 11
0
0 0 880 0
1 1
-4 -14 3 -6
2 R9
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
961 0 0
2
45174.3 4
0
9 Resistor~
219 421 442 0 2 5
0 11 8
0
0 0 880 90
1 5
11 0 18 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3178 0 0
2
45174.3 3
0
9 Resistor~
219 518 443 0 2 5
0 11 8
0
0 0 880 90
2 14
8 0 22 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3409 0 0
2
45174.3 1
0
9 Resistor~
219 518 311 0 2 5
0 15 16
0
0 0 880 90
2 12
8 0 22 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3951 0 0
2
45174.3 0
0
9 Resistor~
219 469 263 0 2 5
0 14 16
0
0 0 880 0
1 2
-4 -14 3 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
8885 0 0
2
45174.3 0
0
9 Resistor~
219 421 310 0 2 5
0 15 14
0
0 0 880 90
1 5
11 0 18 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3780 0 0
2
45174.3 0
0
9 Resistor~
219 384 356 0 2 5
0 12 15
0
0 0 880 0
1 1
-4 -14 3 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9265 0 0
2
45174.3 0
0
9 Resistor~
219 382 263 0 2 5
0 13 14
0
0 0 880 0
1 3
-4 -14 3 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9442 0 0
2
45174.3 0
0
19
2 4 2 0 0 16528 0 6 1 0 0 5
421 668
421 639
356 639
356 657
279 657
1 1 3 0 0 4224 0 1 6 0 0 5
279 707
358 707
358 732
421 732
421 704
2 2 4 0 0 4224 0 7 9 0 0 3
421 547
421 518
400 518
1 1 5 0 0 4224 0 2 8 0 0 4
279 586
358 586
358 611
366 611
4 1 6 0 0 4224 0 2 9 0 0 4
279 536
356 536
356 518
364 518
2 1 7 0 0 8320 0 8 7 0 0 3
402 611
421 611
421 583
2 0 8 0 0 4096 0 12 0 0 12 2
421 424
421 395
1 1 9 0 0 4224 0 3 11 0 0 4
279 463
358 463
358 488
366 488
4 1 10 0 0 4224 0 3 10 0 0 4
279 413
356 413
356 395
364 395
0 1 11 0 0 4096 0 0 12 11 0 2
421 488
421 460
1 2 11 0 0 8320 0 13 11 0 0 3
518 461
518 488
402 488
2 2 8 0 0 4224 0 10 13 0 0 3
400 395
518 395
518 425
1 1 12 0 0 4224 0 5 17 0 0 4
279 331
358 331
358 356
366 356
4 1 13 0 0 4224 0 5 18 0 0 4
279 281
356 281
356 263
364 263
2 0 14 0 0 4096 0 16 0 0 19 2
421 292
421 263
0 1 15 0 0 4096 0 0 16 17 0 2
421 356
421 328
1 2 15 0 0 8320 0 14 17 0 0 3
518 329
518 356
402 356
2 2 16 0 0 4224 0 15 14 0 0 3
487 263
518 263
518 293
2 1 14 0 0 4224 0 18 15 0 0 2
400 263
451 263
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
