CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
120 0 30 150 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
50 C:\Users\Edu\AppData\Local\Temp\IXP001.TMP\BOM.DAT
0 7
5 4 0.500000 0.500000
176 80 1534 803
9437202 0
0
6 Title:
5 Name:
0
0
0
40
13 Logic Switch~
5 206 185 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
6 Enable
-20 -26 22 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3674 0 0
2
45219.3 0
0
13 Logic Switch~
5 205 301 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5697 0 0
2
45219.3 2
0
13 Logic Switch~
5 204 371 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3805 0 0
2
45219.3 1
0
13 Logic Switch~
5 205 334 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5219 0 0
2
45219.3 0
0
13 Logic Switch~
5 204 242 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
6 Enable
-20 -26 22 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3795 0 0
2
45219.3 0
0
5 4049~
219 300 415 0 2 22
0 4 3
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
3637 0 0
2
45219.3 0
0
5 4049~
219 479 491 0 2 22
0 27 11
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
3226 0 0
2
45219.3 3
0
5 4049~
219 479 556 0 2 22
0 25 9
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
6966 0 0
2
45219.3 2
0
5 4049~
219 478 524 0 2 22
0 26 10
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
9796 0 0
2
45219.3 1
0
5 4049~
219 480 586 0 2 22
0 24 8
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
5952 0 0
2
45219.3 0
0
7 74LS138
19 373 398 0 14 29
0 7 6 5 3 2 2 31 30 29
28 27 26 25 24
0
0 0 5104 0
7 74LS138
-25 -61 24 -53
2 U4
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 0 0 0 0
1 U
3649 0 0
2
45219.3 0
0
5 4049~
219 476 393 0 2 22
0 30 14
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 2 0
1 U
3716 0 0
2
45219.3 2
0
5 4049~
219 478 455 0 2 22
0 28 12
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 2 0
1 U
4797 0 0
2
45219.3 1
0
5 4049~
219 477 425 0 2 22
0 29 13
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 2 0
1 U
4681 0 0
2
45219.3 0
0
5 4049~
219 465 86 0 2 22
0 39 23
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
9730 0 0
2
45219.3 8
0
5 4049~
219 466 124 0 2 22
0 38 22
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 1 0
1 U
9874 0 0
2
45219.3 7
0
5 4049~
219 468 160 0 2 22
0 37 21
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 1 0
1 U
364 0 0
2
45219.3 6
0
5 4049~
219 472 263 0 2 22
0 34 18
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 1 0
1 U
3656 0 0
2
45219.3 5
0
5 4049~
219 470 229 0 2 22
0 35 19
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 1 0
1 U
3131 0 0
2
45219.3 4
0
5 4049~
219 477 360 0 2 22
0 31 15
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 2 0
1 U
6772 0 0
2
45219.3 3
0
5 4049~
219 474 329 0 2 22
0 32 16
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 2 0
1 U
9557 0 0
2
45219.3 2
0
5 4049~
219 473 295 0 2 22
0 33 17
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 2 0
1 U
5789 0 0
2
45219.3 1
0
5 4049~
219 469 192 0 2 22
0 36 20
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 1 0
1 U
7328 0 0
2
45219.3 0
0
14 Logic Display~
6 892 40 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4799 0 0
2
45219.3 15
0
14 Logic Display~
6 712 40 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9196 0 0
2
45219.3 14
0
14 Logic Display~
6 734 40 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3857 0 0
2
45219.3 13
0
14 Logic Display~
6 670 40 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7125 0 0
2
45219.3 12
0
14 Logic Display~
6 690 40 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3641 0 0
2
45219.3 11
0
14 Logic Display~
6 757 40 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9821 0 0
2
45219.3 10
0
14 Logic Display~
6 823 40 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3187 0 0
2
45219.3 9
0
14 Logic Display~
6 778 40 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
762 0 0
2
45219.3 8
0
14 Logic Display~
6 800 40 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
39 0 0
2
45219.3 7
0
14 Logic Display~
6 846 40 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9450 0 0
2
45219.3 6
0
14 Logic Display~
6 869 40 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3236 0 0
2
45219.3 5
0
14 Logic Display~
6 624 40 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3321 0 0
2
45219.3 4
0
14 Logic Display~
6 602 40 0 1 2
10 21
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8879 0 0
2
45219.3 3
0
14 Logic Display~
6 581 40 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5433 0 0
2
45219.3 2
0
14 Logic Display~
6 559 40 0 1 2
10 23
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3679 0 0
2
45219.3 1
0
14 Logic Display~
6 648 40 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9342 0 0
2
45219.3 0
0
7 74LS138
19 371 274 0 14 29
0 7 6 5 4 2 2 39 38 37
36 35 34 33 32
0
0 0 5104 0
7 74LS138
-25 -61 24 -53
2 U1
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 0 0 0 0
1 U
3623 0 0
2
45219.3 0
0
45
0 0 2 0 0 4224 0 0 0 2 4 3
246 185
246 429
335 429
1 0 2 0 0 16 0 1 0 0 3 3
218 185
333 185
333 305
6 5 2 0 0 0 0 40 40 0 0 2
333 310
333 301
5 6 2 0 0 0 0 11 11 0 0 2
335 425
335 434
2 4 3 0 0 12416 0 6 11 0 0 4
321 415
327 415
327 416
341 416
0 1 4 0 0 4224 0 0 6 7 0 2
285 242
285 415
1 4 4 0 0 0 0 5 40 0 0 4
216 242
325 242
325 292
339 292
0 3 5 0 0 8192 0 0 11 9 0 3
297 371
297 389
341 389
1 3 5 0 0 8320 0 3 40 0 0 4
216 371
297 371
297 265
339 265
0 2 6 0 0 4096 0 0 11 11 0 3
312 334
312 380
341 380
1 2 6 0 0 4224 0 4 40 0 0 4
217 334
312 334
312 256
339 256
0 1 7 0 0 4096 0 0 11 13 0 3
319 301
319 371
341 371
1 1 7 0 0 4224 0 2 40 0 0 4
217 301
319 301
319 247
339 247
1 2 8 0 0 4224 0 24 10 0 0 3
892 58
892 586
501 586
1 2 9 0 0 4224 0 34 8 0 0 3
869 58
869 556
500 556
1 2 10 0 0 4224 0 33 9 0 0 3
846 58
846 524
499 524
1 2 11 0 0 4224 0 30 7 0 0 3
823 58
823 491
500 491
1 2 12 0 0 4224 0 32 13 0 0 3
800 58
800 455
499 455
1 2 13 0 0 4224 0 31 14 0 0 3
778 58
778 425
498 425
2 1 14 0 0 8320 0 12 29 0 0 3
497 393
757 393
757 58
2 1 15 0 0 8320 0 20 26 0 0 3
498 360
734 360
734 58
2 1 16 0 0 8320 0 21 25 0 0 3
495 329
712 329
712 58
2 1 17 0 0 8320 0 22 28 0 0 3
494 295
690 295
690 58
2 1 18 0 0 8320 0 18 27 0 0 3
493 263
670 263
670 58
2 1 19 0 0 8320 0 19 39 0 0 3
491 229
648 229
648 58
2 1 20 0 0 4224 0 23 35 0 0 3
490 192
624 192
624 58
2 1 21 0 0 4224 0 17 36 0 0 3
489 160
602 160
602 58
2 1 22 0 0 4224 0 16 37 0 0 3
487 124
581 124
581 58
2 1 23 0 0 4224 0 15 38 0 0 3
486 86
559 86
559 58
14 1 24 0 0 8320 0 11 10 0 0 4
411 434
422 434
422 586
465 586
13 1 25 0 0 8320 0 11 8 0 0 4
411 425
428 425
428 556
464 556
12 1 26 0 0 8320 0 11 9 0 0 4
411 416
433 416
433 524
463 524
11 1 27 0 0 8320 0 11 7 0 0 4
411 407
440 407
440 491
464 491
10 1 28 0 0 8320 0 11 13 0 0 4
411 398
445 398
445 455
463 455
9 1 29 0 0 4224 0 11 14 0 0 4
411 389
449 389
449 425
462 425
8 1 30 0 0 4224 0 11 12 0 0 4
411 380
453 380
453 393
461 393
7 1 31 0 0 4224 0 11 20 0 0 4
411 371
453 371
453 360
462 360
14 1 32 0 0 4224 0 40 21 0 0 4
409 310
451 310
451 329
459 329
13 1 33 0 0 4224 0 40 22 0 0 4
409 301
450 301
450 295
458 295
12 1 34 0 0 4224 0 40 18 0 0 4
409 292
449 292
449 263
457 263
11 1 35 0 0 8320 0 40 19 0 0 4
409 283
442 283
442 229
455 229
10 1 36 0 0 8320 0 40 23 0 0 4
409 274
436 274
436 192
454 192
9 1 37 0 0 8320 0 40 17 0 0 4
409 265
427 265
427 160
453 160
8 1 38 0 0 8320 0 40 16 0 0 4
409 256
422 256
422 124
451 124
7 1 39 0 0 8320 0 40 15 0 0 4
409 247
416 247
416 86
450 86
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
