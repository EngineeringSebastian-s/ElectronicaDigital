CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
160 140 30 200 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
50 C:\Users\Edu\AppData\Local\Temp\IXP000.TMP\BOM.DAT
0 7
2 4 0.499308 0.500000
344 176 1702 537
9961490 0
0
6 Title:
5 Name:
0
0
0
7
8 Battery~
219 219 349 0 2 5
0 3 2
0
0 0 880 0
3 10V
12 -2 33 6
2 V1
16 -12 30 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
7361 0 0
2
45177.9 0
0
11 Multimeter~
205 221 230 0 21 21
0 3 7 8 4 0 0 0 0 0
32 50 52 46 54 57 109 65 0 0
0 86
0
0 0 16464 0
6 1.000u
-21 -19 21 -11
3 MM0
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
4747 0 0
2
45177.9 0
0
7 Ground~
168 616 380 0 1 3
0 9
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 0 0 0 0
3 GND
972 0 0
2
45177.9 0
0
9 Resistor~
219 479 335 0 2 5
0 5 6
0
0 0 880 90
3 350
5 0 26 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3472 0 0
2
45177.9 0
0
9 Resistor~
219 407 332 0 2 5
0 5 6
0
0 0 880 90
3 150
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9998 0 0
2
45177.9 0
0
9 Resistor~
219 353 375 0 2 5
0 2 5
0
0 0 880 0
3 200
-10 -14 11 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3536 0 0
2
45177.9 0
0
9 Resistor~
219 353 288 0 2 5
0 4 6
0
0 0 880 0
3 100
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
4597 0 0
2
45177.9 0
0
7
2 1 2 0 0 8320 0 1 6 0 0 3
219 360
219 375
335 375
1 1 3 0 0 4224 0 2 1 0 0 4
196 253
196 321
219 321
219 336
4 1 4 0 0 8320 0 2 7 0 0 3
246 253
246 288
335 288
0 1 5 0 0 4224 0 0 4 7 0 3
407 375
479 375
479 353
0 2 6 0 0 4240 0 0 4 6 0 3
407 288
479 288
479 317
2 2 6 0 0 0 0 7 5 0 0 3
371 288
407 288
407 314
2 1 5 0 0 0 0 6 5 0 0 3
371 375
407 375
407 350
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
