CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
160 10 30 150 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
50 C:\Users\Edu\AppData\Local\Temp\IXP000.TMP\BOM.DAT
0 7
2 4 0.323651 0.500000
344 176 1702 410
9961490 0
0
6 Title:
5 Name:
0
0
0
18
8 Battery~
219 407 278 0 2 5
0 3 4
0
0 0 880 90
3 12v
-11 -21 10 -13
2 V1
-7 -31 7 -23
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
5130 0 0
2
45172.6 0
0
7 Ground~
168 685 375 0 1 3
0 11
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 0 0 0 0
3 GND
391 0 0
2
45172.6 0
0
11 Multimeter~
205 348 254 0 21 21
0 3 12 13 2 0 0 0 0 0
32 50 46 50 52 57 32 65 0 0
0 86
0
0 0 16464 90
6 1.000u
-21 -19 21 -11
3 MM0
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 0 0 0 0
1 V
3124 0 0
2
45172.6 0
0
9 Resistor~
219 605 222 0 2 5
0 7 6
0
0 0 880 0
1 2
-4 -14 3 -6
3 R15
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3421 0 0
2
45172.6 0
0
9 Resistor~
219 503 221 0 2 5
0 2 7
0
0 0 880 0
1 6
-4 -14 3 -6
3 R14
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
8157 0 0
2
45172.6 0
0
9 Resistor~
219 363 221 0 2 5
0 8 2
0
0 0 880 0
2 12
-7 -14 7 -6
3 R13
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
5572 0 0
2
45172.6 0
0
9 Resistor~
219 651 254 0 2 5
0 5 6
0
0 0 880 90
1 5
11 0 18 8
3 R12
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
8901 0 0
2
45172.6 0
0
9 Resistor~
219 559 250 0 2 5
0 5 7
0
0 0 880 90
2 10
8 0 22 8
3 R11
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7361 0 0
2
45172.6 0
0
9 Resistor~
219 303 258 0 2 5
0 4 8
0
0 0 880 90
2 12
8 0 22 8
3 R10
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
4747 0 0
2
45172.6 0
0
9 Resistor~
219 210 257 0 2 5
0 9 8
0
0 0 880 90
1 7
11 0 18 8
2 R9
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
972 0 0
2
45172.6 0
0
9 Resistor~
219 501 295 0 2 5
0 4 5
0
0 0 880 0
1 4
-4 -14 3 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3472 0 0
2
45172.6 0
0
9 Resistor~
219 262 295 0 2 5
0 9 4
0
0 0 880 0
2 10
-7 -14 7 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9998 0 0
2
45172.6 0
0
9 Resistor~
219 558 366 0 2 5
0 4 5
0
0 0 880 0
2 10
-7 -14 7 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3536 0 0
2
45172.6 0
0
9 Resistor~
219 309 367 0 2 5
0 9 4
0
0 0 880 0
2 10
-7 -14 7 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
4597 0 0
2
45172.6 0
0
9 Resistor~
219 603 185 0 2 5
0 7 6
0
0 0 880 0
1 2
-4 -14 3 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3835 0 0
2
45172.6 0
0
9 Resistor~
219 504 185 0 2 5
0 2 7
0
0 0 880 0
1 6
-4 -14 3 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3670 0 0
2
45172.6 0
0
9 Resistor~
219 365 185 0 2 5
0 10 2
0
0 0 880 0
1 8
-4 -14 3 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
5616 0 0
2
45172.6 0
0
9 Resistor~
219 261 185 0 2 5
0 8 10
0
0 0 880 0
1 4
-4 -14 3 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9323 0 0
2
45172.6 0
0
25
4 0 2 0 0 4112 0 3 0 0 5 4
365 235
425 235
425 221
426 221
1 1 3 0 0 4224 0 1 3 0 0 4
397 275
372 275
372 285
365 285
2 0 4 0 0 8192 0 1 0 0 4 4
421 275
434 275
434 295
427 295
0 0 4 0 0 4096 0 0 0 15 22 2
427 295
427 367
0 0 2 0 0 0 0 0 0 24 10 2
426 185
426 221
1 0 5 0 0 4096 0 8 0 0 14 2
559 268
559 295
2 0 6 0 0 4096 0 4 0 0 18 2
623 222
651 222
0 1 7 0 0 8192 0 0 4 9 0 3
558 221
558 222
587 222
2 0 7 0 0 4096 0 5 0 0 17 2
521 221
559 221
2 1 2 0 0 4224 0 6 5 0 0 2
381 221
485 221
0 1 8 0 0 4096 0 0 6 13 0 2
303 221
345 221
1 0 4 0 0 0 0 9 0 0 15 2
303 276
303 295
0 2 8 0 0 4224 0 0 9 21 0 3
210 221
303 221
303 240
2 0 5 0 0 4224 0 11 0 0 19 2
519 295
651 295
2 1 4 0 0 4224 0 12 11 0 0 2
280 295
483 295
0 1 9 0 0 4096 0 0 12 20 0 2
210 295
244 295
0 2 7 0 0 4096 0 0 8 23 0 2
559 185
559 232
2 2 6 0 0 8320 0 15 7 0 0 3
621 185
651 185
651 236
2 1 5 0 0 0 0 13 7 0 0 3
576 366
651 366
651 272
1 1 9 0 0 4224 0 10 14 0 0 3
210 275
210 367
291 367
1 2 8 0 0 0 0 18 10 0 0 3
243 185
210 185
210 239
2 1 4 0 0 128 0 14 13 0 0 4
327 367
525 367
525 366
540 366
2 1 7 0 0 4224 0 16 15 0 0 2
522 185
585 185
2 1 2 0 0 0 0 17 16 0 0 2
383 185
486 185
2 1 10 0 0 4224 0 18 17 0 0 2
279 185
347 185
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
