CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
50 C:\Users\Edu\AppData\Local\Temp\IXP001.TMP\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
49
13 Logic Switch~
5 223 681 0 1 11
0 8
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 C1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7168 0 0
2
45198.6 3
0
13 Logic Switch~
5 187 683 0 1 11
0 4
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 B1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
631 0 0
2
45198.6 2
0
13 Logic Switch~
5 148 683 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9466 0 0
2
45198.6 1
0
13 Logic Switch~
5 262 681 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 D1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3266 0 0
2
45198.6 0
0
13 Logic Switch~
5 263 117 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 D
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7693 0 0
2
45198.6 0
0
13 Logic Switch~
5 149 119 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3723 0 0
2
45198.6 1
0
13 Logic Switch~
5 188 119 0 1 11
0 30
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3440 0 0
2
45198.6 2
0
13 Logic Switch~
5 224 117 0 1 11
0 27
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 C
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6263 0 0
2
45198.6 3
0
8 3-In OR~
219 757 1040 0 4 22
0 12 14 13 11
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 8 0
1 U
4900 0 0
2
45198.6 0
0
8 4-In OR~
219 653 885 0 5 22
0 18 17 2 15 12
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U11A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 12 0
1 U
8783 0 0
2
45198.6 0
0
5 4073~
219 448 1116 0 4 22
0 20 8 19 13
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U10C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 11 0
1 U
3221 0 0
2
45198.6 0
0
5 4073~
219 445 1041 0 4 22
0 22 8 21 14
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U10B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 11 0
1 U
3215 0 0
2
45198.6 0
0
5 4073~
219 442 979 0 4 22
0 10 4 9 15
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U10A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 11 0
1 U
7903 0 0
2
45198.6 0
0
5 4073~
219 441 917 0 4 22
0 10 4 5 2
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 10 0
1 U
7121 0 0
2
45198.6 0
0
5 4073~
219 435 846 0 4 22
0 10 23 9 17
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 10 0
1 U
4484 0 0
2
45198.6 0
0
5 4073~
219 436 780 0 4 22
0 4 24 8 18
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 10 0
1 U
5996 0 0
2
45198.6 0
0
5 4049~
219 317 771 0 2 22
0 8 24
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 9 0
1 U
7804 0 0
2
45198.6 16
0
5 4049~
219 320 847 0 2 22
0 8 23
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 9 0
1 U
5523 0 0
2
45198.6 15
0
5 4049~
219 324 938 0 2 22
0 8 5
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 5 0
1 U
3330 0 0
2
45198.6 14
0
5 4049~
219 327 1022 0 2 22
0 4 22
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 5 0
1 U
3465 0 0
2
45198.6 13
0
5 4049~
219 328 1066 0 2 22
0 9 21
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 5 0
1 U
8396 0 0
2
45198.6 12
0
5 4049~
219 332 1099 0 2 22
0 10 20
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 5 0
1 U
3685 0 0
2
45198.6 11
0
5 4049~
219 336 1150 0 2 22
0 9 19
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 5 0
1 U
7849 0 0
2
45198.6 10
0
14 Logic Display~
6 881 818 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6343 0 0
2
45198.6 4
0
14 Logic Display~
6 882 254 0 1 2
10 32
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7376 0 0
2
45198.6 4
0
5 4071~
219 797 359 0 3 22
0 33 34 32
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
9156 0 0
2
45198.6 5
0
5 4071~
219 602 537 0 3 22
0 36 35 34
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U5D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 6 0
1 U
5776 0 0
2
45198.6 6
0
5 4071~
219 690 314 0 3 22
0 40 39 33
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 6 0
1 U
7207 0 0
2
45198.6 7
0
5 4071~
219 600 396 0 3 22
0 38 37 39
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
4459 0 0
2
45198.6 8
0
5 4071~
219 594 249 0 3 22
0 42 41 40
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
3760 0 0
2
45198.6 9
0
5 4049~
219 337 586 0 2 22
0 28 44
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 5 0
1 U
754 0 0
2
45198.6 10
0
5 4049~
219 333 535 0 2 22
0 31 45
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 4 0
1 U
9767 0 0
2
45198.6 11
0
5 4049~
219 329 502 0 2 22
0 28 47
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 4 0
1 U
7978 0 0
2
45198.6 12
0
5 4049~
219 328 458 0 2 22
0 30 48
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 4 0
1 U
3142 0 0
2
45198.6 13
0
5 4049~
219 325 374 0 2 22
0 27 52
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 4 0
1 U
3284 0 0
2
45198.6 14
0
5 4049~
219 321 283 0 2 22
0 27 53
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 4 0
1 U
659 0 0
2
45198.6 15
0
5 4049~
219 318 207 0 2 22
0 27 54
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 4 0
1 U
3800 0 0
2
45198.6 16
0
5 4081~
219 409 197 0 3 22
0 30 54 49
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
6792 0 0
2
45198.6 17
0
5 4081~
219 411 269 0 3 22
0 31 53 50
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
3701 0 0
2
45198.6 18
0
5 4081~
219 413 338 0 3 22
0 31 30 51
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
6316 0 0
2
45198.6 19
0
5 4081~
219 415 405 0 3 22
0 31 30 29
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
8734 0 0
2
45198.6 20
0
5 4081~
219 416 471 0 3 22
0 48 27 46
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1E
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
7988 0 0
2
45198.6 21
0
5 4081~
219 418 542 0 3 22
0 45 27 43
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1F
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
3217 0 0
2
45198.6 22
0
5 4081~
219 479 216 0 3 22
0 49 27 42
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
3965 0 0
2
45198.6 23
0
5 4081~
219 479 291 0 3 22
0 50 28 41
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
8239 0 0
2
45198.6 24
0
5 4081~
219 482 367 0 3 22
0 51 52 38
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
828 0 0
2
45198.6 25
0
5 4081~
219 484 434 0 3 22
0 29 28 37
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
6187 0 0
2
45198.6 26
0
5 4081~
219 485 506 0 3 22
0 46 47 36
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
7107 0 0
2
45198.6 27
0
5 4081~
219 486 575 0 3 22
0 43 44 35
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 3 0
1 U
6433 0 0
2
45198.6 28
0
83
3 4 2 0 0 12416 0 10 14 0 0 4
636 890
578 890
578 917
462 917
0 0 3 0 0 4224 0 0 0 0 0 2
579 882
578 882
0 2 4 0 0 12288 0 0 14 37 0 4
187 923
202 923
202 917
417 917
2 3 5 0 0 4224 0 19 14 0 0 4
345 938
404 938
404 926
417 926
0 0 6 0 0 0 0 0 0 0 0 2
187 1120
187 1120
0 0 7 0 0 0 0 0 0 0 0 2
148 1122
148 1122
0 2 8 0 0 4096 0 0 11 36 0 3
223 1115
424 1115
424 1116
0 1 9 0 0 12288 0 0 21 35 0 4
262 1064
277 1064
277 1066
313 1066
0 2 8 0 0 0 0 0 12 36 0 4
223 1044
238 1044
238 1041
421 1041
0 3 9 0 0 4096 0 0 13 35 0 3
262 1000
418 1000
418 988
0 2 4 0 0 12288 0 0 13 37 0 4
187 978
202 978
202 979
418 979
0 1 10 0 0 4096 0 0 13 38 0 3
148 960
418 960
418 970
0 1 8 0 0 0 0 0 19 36 0 2
223 938
309 938
0 1 10 0 0 0 0 0 14 38 0 4
148 893
388 893
388 908
417 908
0 3 9 0 0 0 0 0 15 35 0 3
262 864
411 864
411 855
0 1 8 0 0 0 0 0 18 36 0 2
223 847
305 847
0 1 10 0 0 0 0 0 15 38 0 3
148 824
411 824
411 837
0 3 8 0 0 0 0 0 16 36 0 2
223 789
412 789
0 1 8 0 0 0 0 0 17 36 0 2
223 771
302 771
0 1 4 0 0 0 0 0 16 37 0 5
187 710
365 710
365 755
412 755
412 771
4 1 11 0 0 8320 0 9 24 0 0 3
790 1040
881 1040
881 836
5 1 12 0 0 8320 0 10 9 0 0 4
686 885
731 885
731 1031
744 1031
4 3 13 0 0 4240 0 11 9 0 0 6
469 1116
603 1116
603 1089
732 1089
732 1049
744 1049
4 2 14 0 0 12416 0 12 9 0 0 4
466 1041
588 1041
588 1040
745 1040
4 4 15 0 0 4224 0 13 10 0 0 5
463 979
578 979
578 964
636 964
636 899
0 0 16 0 0 4224 0 0 0 0 0 2
579 831
578 831
4 2 17 0 0 4224 0 15 10 0 0 4
456 846
572 846
572 881
636 881
4 1 18 0 0 4224 0 16 10 0 0 5
457 780
572 780
572 832
636 832
636 872
2 3 19 0 0 4224 0 23 11 0 0 4
357 1150
398 1150
398 1125
424 1125
2 1 20 0 0 12416 0 22 11 0 0 4
353 1099
368 1099
368 1107
424 1107
2 3 21 0 0 4224 0 21 12 0 0 4
349 1066
396 1066
396 1050
421 1050
2 1 22 0 0 12416 0 20 12 0 0 4
348 1022
383 1022
383 1032
421 1032
2 2 23 0 0 4224 0 18 15 0 0 3
341 847
411 847
411 846
2 2 24 0 0 4224 0 17 16 0 0 5
338 771
376 771
376 778
412 778
412 780
1 1 9 0 0 8320 0 23 4 0 0 3
321 1150
262 1150
262 693
1 0 8 0 0 4224 0 1 0 0 0 2
223 693
223 1117
1 1 4 0 0 4224 0 2 20 0 0 3
187 695
187 1022
312 1022
1 1 10 0 0 4224 0 3 22 0 0 3
148 695
148 1099
317 1099
0 0 25 0 0 0 0 0 0 0 0 2
188 556
188 556
0 0 26 0 0 0 0 0 0 0 0 2
149 558
149 558
0 2 27 0 0 4096 0 0 43 81 0 2
224 551
394 551
0 1 28 0 0 12288 0 0 33 80 0 4
263 500
278 500
278 502
314 502
0 2 27 0 0 0 0 0 42 81 0 2
224 480
392 480
3 1 29 0 0 8320 0 41 47 0 0 4
436 405
452 405
452 425
460 425
0 2 28 0 0 4096 0 0 47 80 0 3
263 436
460 436
460 443
0 2 30 0 0 4096 0 0 41 82 0 2
188 414
391 414
0 1 31 0 0 4096 0 0 41 83 0 2
149 396
391 396
0 1 27 0 0 0 0 0 35 81 0 2
224 374
310 374
0 2 30 0 0 0 0 0 40 82 0 2
188 347
389 347
0 1 31 0 0 0 0 0 40 83 0 2
149 329
389 329
0 2 28 0 0 0 0 0 45 80 0 2
263 300
455 300
0 1 27 0 0 0 0 0 36 81 0 2
224 283
306 283
0 1 31 0 0 0 0 0 39 83 0 2
149 260
387 260
0 2 27 0 0 4096 0 0 44 81 0 2
224 225
455 225
0 1 27 0 0 0 0 0 37 81 0 2
224 207
303 207
0 1 30 0 0 0 0 0 38 82 0 4
188 146
366 146
366 188
385 188
3 1 32 0 0 8320 0 26 25 0 0 3
830 359
882 359
882 272
3 1 33 0 0 12416 0 28 26 0 0 4
723 314
732 314
732 350
784 350
3 2 34 0 0 8320 0 27 26 0 0 4
635 537
710 537
710 368
784 368
3 2 35 0 0 4224 0 49 27 0 0 4
507 575
581 575
581 546
589 546
3 1 36 0 0 4224 0 48 27 0 0 4
506 506
581 506
581 528
589 528
3 2 37 0 0 4224 0 47 29 0 0 4
505 434
579 434
579 405
587 405
3 1 38 0 0 4224 0 46 29 0 0 4
503 367
579 367
579 387
587 387
3 2 39 0 0 8320 0 29 28 0 0 4
633 396
669 396
669 323
677 323
3 1 40 0 0 8320 0 30 28 0 0 4
627 249
669 249
669 305
677 305
3 2 41 0 0 4224 0 45 30 0 0 4
500 291
573 291
573 258
581 258
3 1 42 0 0 4224 0 44 30 0 0 4
500 216
573 216
573 240
581 240
3 1 43 0 0 8320 0 43 49 0 0 4
439 542
454 542
454 566
462 566
2 2 44 0 0 4224 0 31 49 0 0 4
358 586
454 586
454 584
462 584
2 1 45 0 0 4224 0 32 43 0 0 4
354 535
386 535
386 533
394 533
3 1 46 0 0 8320 0 42 48 0 0 4
437 471
448 471
448 497
461 497
2 2 47 0 0 4224 0 33 48 0 0 4
350 502
437 502
437 515
461 515
2 1 48 0 0 4224 0 34 42 0 0 4
349 458
384 458
384 462
392 462
3 1 49 0 0 4224 0 38 44 0 0 4
430 197
447 197
447 207
455 207
3 1 50 0 0 4224 0 39 45 0 0 4
432 269
447 269
447 282
455 282
3 1 51 0 0 8320 0 40 46 0 0 4
434 338
450 338
450 358
458 358
2 2 52 0 0 4224 0 35 46 0 0 4
346 374
450 374
450 376
458 376
2 2 53 0 0 4224 0 36 39 0 0 4
342 283
379 283
379 278
387 278
2 2 54 0 0 4224 0 37 38 0 0 4
339 207
377 207
377 206
385 206
1 1 28 0 0 8320 0 31 5 0 0 3
322 586
263 586
263 129
1 0 27 0 0 4224 0 8 0 0 0 2
224 129
224 553
1 1 30 0 0 4224 0 7 34 0 0 3
188 131
188 458
313 458
1 1 31 0 0 4224 0 6 32 0 0 3
149 131
149 535
318 535
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
