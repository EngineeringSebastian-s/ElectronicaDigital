CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
120 110 30 150 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
50 C:\Users\Edu\AppData\Local\Temp\IXP000.TMP\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1702 537
9961490 0
0
6 Title:
5 Name:
0
0
0
23
7 Ground~
168 941 214 0 1 3
0 15
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 0 0 0 0
3 GND
6369 0 0
2
45177.9 0
0
11 Multimeter~
205 212 343 0 21 21
0 7 16 17 9 0 0 0 0 0
32 51 57 52 46 55 32 32 0 0
4 73
0
0 0 16464 90
6 1.000u
-21 -19 21 -11
3 MM0
-11 -29 10 -21
0
0
31 R1%D %1 %2 1E-9
%D %4 %2 DC %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
73 0 0 0 1 0 0 0
1 I
9172 0 0
2
45177.9 6
0
9 Resistor~
219 932 362 0 2 5
0 3 4
0
0 0 880 90
3 530
8 0 29 8
3 R21
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7100 0 0
2
45177.9 90
0
9 Resistor~
219 557 277 0 2 5
0 5 6
0
0 0 880 90
3 900
8 0 29 8
3 R20
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3820 0 0
2
45177.9 91
0
9 Resistor~
219 421 415 0 2 5
0 5 6
0
0 0 880 90
3 500
8 0 29 8
3 R19
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7678 0 0
2
45177.9 92
0
9 Resistor~
219 317 294 0 2 5
0 7 10
0
0 0 880 90
3 200
8 0 29 8
3 R18
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
961 0 0
2
45177.9 93
0
9 Resistor~
219 817 470 0 2 5
0 8 3
0
0 0 880 0
4 3.5k
-14 -14 14 -6
3 R17
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3178 0 0
2
45177.9 94
0
9 Resistor~
219 866 407 0 2 5
0 3 11
0
0 0 880 90
3 150
8 0 29 8
3 R16
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3409 0 0
2
45177.9 95
0
9 Resistor~
219 865 293 0 2 5
0 11 4
0
0 0 880 90
3 280
8 0 29 8
3 R15
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3951 0 0
2
45177.9 96
0
9 Resistor~
219 803 233 0 2 5
0 2 4
0
0 0 880 0
3 380
-10 -14 11 -6
3 R14
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8885 0 0
2
45177.9 97
0
9 Resistor~
219 669 407 0 2 5
0 8 2
0
0 0 880 90
2 4k
11 0 25 8
3 R13
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3780 0 0
2
45177.9 98
0
9 Resistor~
219 729 409 0 2 5
0 8 12
0
0 0 880 90
3 400
8 0 29 8
3 R12
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9265 0 0
2
45177.9 99
0
9 Resistor~
219 729 306 0 2 5
0 12 2
0
0 0 880 90
3 520
8 0 29 8
3 R11
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9442 0 0
2
45177.9 100
0
9 Resistor~
219 616 470 0 2 5
0 5 8
0
0 0 880 0
3 350
-10 -14 11 -6
3 R10
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9424 0 0
2
45177.9 101
0
9 Resistor~
219 613 351 0 2 5
0 5 2
0
0 0 880 0
3 600
-10 -14 11 -6
2 R9
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9968 0 0
2
45177.9 102
0
9 Resistor~
219 614 233 0 2 5
0 6 2
0
0 0 880 0
4 2.1k
-14 -14 14 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9281 0 0
2
45177.9 103
0
9 Resistor~
219 497 419 0 2 5
0 5 13
0
0 0 880 90
4 850k
2 0 30 8
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8464 0 0
2
45177.9 104
0
9 Resistor~
219 497 357 0 2 5
0 13 14
0
0 0 880 90
3 850
5 0 26 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7168 0 0
2
45177.9 105
0
9 Resistor~
219 497 295 0 2 5
0 14 6
0
0 0 880 90
3 750
5 0 26 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3171 0 0
2
45177.9 106
0
9 Resistor~
219 374 470 0 2 5
0 7 5
0
0 0 880 0
3 100
-10 -14 11 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4139 0 0
2
45177.9 107
0
9 Resistor~
219 372 352 0 2 5
0 7 6
0
0 0 880 0
4 300k
-14 -14 14 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6435 0 0
2
45177.9 108
0
9 Resistor~
219 367 233 0 2 5
0 6 10
0
0 0 880 180
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5283 0 0
2
45177.9 109
0
9 Resistor~
219 248 267 0 2 5
0 10 9
0
0 0 880 270
3 220
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6874 0 0
2
45177.9 110
0
31
2 0 2 0 0 4096 0 15 0 0 2 2
631 351
669 351
2 0 2 0 0 4224 0 11 0 0 4 2
669 389
669 233
2 0 2 0 0 0 0 13 0 0 4 2
729 288
729 233
2 1 2 0 0 0 0 16 10 0 0 2
632 233
785 233
0 1 3 0 0 4224 0 0 3 20 0 3
866 440
932 440
932 380
0 2 4 0 0 8320 0 0 3 22 0 3
865 271
932 271
932 344
1 0 5 0 0 4096 0 4 0 0 15 2
557 295
557 352
0 2 6 0 0 4096 0 0 4 27 0 2
557 233
557 259
2 0 6 0 0 4096 0 21 0 0 11 2
390 352
421 352
1 0 5 0 0 0 0 5 0 0 24 2
421 433
421 470
0 2 6 0 0 4224 0 0 5 28 0 2
421 233
421 397
0 1 7 0 0 4096 0 0 21 13 0 2
317 352
354 352
1 0 7 0 0 4224 0 6 0 0 14 2
317 312
317 470
1 1 7 0 0 128 0 2 20 0 0 4
229 374
248 374
248 470
356 470
1 0 5 0 0 8192 0 15 0 0 23 3
595 351
557 351
557 470
1 0 8 0 0 4096 0 11 0 0 25 2
669 425
669 470
2 4 9 0 0 4224 0 23 2 0 0 3
248 285
248 324
229 324
0 2 10 0 0 4096 0 0 6 29 0 2
317 233
317 276
1 0 8 0 0 4096 0 7 0 0 25 4
799 470
852 470
852 470
837 470
1 2 3 0 0 0 0 8 7 0 0 3
866 425
866 470
835 470
1 2 11 0 0 4224 0 9 8 0 0 4
865 311
865 372
866 372
866 389
2 2 4 0 0 16 0 10 9 0 0 3
821 233
865 233
865 275
0 1 5 0 0 128 0 0 14 24 0 2
519 470
598 470
2 1 5 0 0 4224 0 20 17 0 0 5
392 470
519 470
519 470
497 470
497 437
2 1 8 0 0 4224 0 14 12 0 0 5
634 470
837 470
837 470
729 470
729 427
2 1 12 0 0 4224 0 12 13 0 0 2
729 391
729 324
0 1 6 0 0 0 0 0 16 28 0 2
518 233
596 233
1 2 6 0 0 0 0 22 19 0 0 5
385 233
518 233
518 233
497 233
497 277
1 2 10 0 0 8320 0 23 22 0 0 3
248 249
248 233
349 233
1 2 13 0 0 4224 0 18 17 0 0 2
497 375
497 401
2 1 14 0 0 4224 0 18 19 0 0 2
497 339
497 313
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
